magic
tech sky130A
magscale 1 2
timestamp 1647800759
<< viali >>
rect 9965 37417 9999 37451
rect 33517 37417 33551 37451
rect 18705 37349 18739 37383
rect 10701 37281 10735 37315
rect 11989 37281 12023 37315
rect 15209 37281 15243 37315
rect 19993 37281 20027 37315
rect 22017 37281 22051 37315
rect 34161 37281 34195 37315
rect 1409 37213 1443 37247
rect 2329 37213 2363 37247
rect 3801 37213 3835 37247
rect 6561 37213 6595 37247
rect 7849 37213 7883 37247
rect 9873 37213 9907 37247
rect 11529 37213 11563 37247
rect 14105 37213 14139 37247
rect 15025 37213 15059 37247
rect 17601 37213 17635 37247
rect 19441 37213 19475 37247
rect 22753 37213 22787 37247
rect 23581 37213 23615 37247
rect 24593 37213 24627 37247
rect 25973 37213 26007 37247
rect 28089 37213 28123 37247
rect 28549 37213 28583 37247
rect 34897 37213 34931 37247
rect 36737 37213 36771 37247
rect 37381 37213 37415 37247
rect 11713 37145 11747 37179
rect 19625 37145 19659 37179
rect 35081 37145 35115 37179
rect 1593 37077 1627 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 22845 37077 22879 37111
rect 24409 37077 24443 37111
rect 27997 37077 28031 37111
rect 37473 37077 37507 37111
rect 10885 36873 10919 36907
rect 19901 36873 19935 36907
rect 20545 36805 20579 36839
rect 22017 36805 22051 36839
rect 24317 36805 24351 36839
rect 27905 36805 27939 36839
rect 35081 36805 35115 36839
rect 1409 36737 1443 36771
rect 2789 36737 2823 36771
rect 3433 36737 3467 36771
rect 10333 36737 10367 36771
rect 10793 36737 10827 36771
rect 13645 36737 13679 36771
rect 17509 36737 17543 36771
rect 19993 36737 20027 36771
rect 20453 36737 20487 36771
rect 21281 36737 21315 36771
rect 21833 36737 21867 36771
rect 24133 36737 24167 36771
rect 33793 36737 33827 36771
rect 34897 36737 34931 36771
rect 36737 36737 36771 36771
rect 37381 36737 37415 36771
rect 3617 36669 3651 36703
rect 4169 36669 4203 36703
rect 12265 36669 12299 36703
rect 13461 36669 13495 36703
rect 17693 36669 17727 36703
rect 18061 36669 18095 36703
rect 22293 36669 22327 36703
rect 24593 36669 24627 36703
rect 27721 36669 27755 36703
rect 29101 36669 29135 36703
rect 1593 36533 1627 36567
rect 2697 36533 2731 36567
rect 21189 36533 21223 36567
rect 34437 36533 34471 36567
rect 37473 36533 37507 36567
rect 3893 36329 3927 36363
rect 12633 36329 12667 36363
rect 17693 36329 17727 36363
rect 19625 36329 19659 36363
rect 35081 36329 35115 36363
rect 1409 36193 1443 36227
rect 3065 36193 3099 36227
rect 3249 36193 3283 36227
rect 10241 36193 10275 36227
rect 12081 36193 12115 36227
rect 21189 36193 21223 36227
rect 22385 36193 22419 36227
rect 22569 36193 22603 36227
rect 25881 36193 25915 36227
rect 26433 36193 26467 36227
rect 36277 36193 36311 36227
rect 36461 36193 36495 36227
rect 38117 36193 38151 36227
rect 3985 36125 4019 36159
rect 12725 36125 12759 36159
rect 17601 36125 17635 36159
rect 24409 36125 24443 36159
rect 25237 36125 25271 36159
rect 34161 36125 34195 36159
rect 34989 36125 35023 36159
rect 35633 36125 35667 36159
rect 11897 36057 11931 36091
rect 25329 36057 25363 36091
rect 26065 36057 26099 36091
rect 35725 35989 35759 36023
rect 11621 35785 11655 35819
rect 36737 35717 36771 35751
rect 11713 35649 11747 35683
rect 23949 35649 23983 35683
rect 34897 35649 34931 35683
rect 38025 35649 38059 35683
rect 24133 35581 24167 35615
rect 24593 35581 24627 35615
rect 35081 35581 35115 35615
rect 37933 35445 37967 35479
rect 24501 35241 24535 35275
rect 35633 35241 35667 35275
rect 36277 35105 36311 35139
rect 36461 35105 36495 35139
rect 38117 35105 38151 35139
rect 1685 35037 1719 35071
rect 24593 35037 24627 35071
rect 35541 35037 35575 35071
rect 1593 34561 1627 34595
rect 37473 34561 37507 34595
rect 1777 34493 1811 34527
rect 2789 34493 2823 34527
rect 37565 34493 37599 34527
rect 36553 34357 36587 34391
rect 2053 34153 2087 34187
rect 36277 34017 36311 34051
rect 36461 34017 36495 34051
rect 38117 34017 38151 34051
rect 2145 33949 2179 33983
rect 26433 33541 26467 33575
rect 38025 33473 38059 33507
rect 24593 33405 24627 33439
rect 24777 33405 24811 33439
rect 37841 33337 37875 33371
rect 18613 33269 18647 33303
rect 36553 33269 36587 33303
rect 24685 33065 24719 33099
rect 19257 32929 19291 32963
rect 19717 32929 19751 32963
rect 36277 32929 36311 32963
rect 19441 32793 19475 32827
rect 36461 32793 36495 32827
rect 38117 32793 38151 32827
rect 19165 32521 19199 32555
rect 24317 32521 24351 32555
rect 36645 32521 36679 32555
rect 19257 32385 19291 32419
rect 24225 32385 24259 32419
rect 36737 32385 36771 32419
rect 37381 32385 37415 32419
rect 1685 32181 1719 32215
rect 36093 32181 36127 32215
rect 37473 32181 37507 32215
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 36277 31841 36311 31875
rect 36461 31841 36495 31875
rect 38117 31841 38151 31875
rect 35817 31773 35851 31807
rect 1593 31705 1627 31739
rect 2053 31433 2087 31467
rect 36553 31365 36587 31399
rect 37381 31365 37415 31399
rect 2145 31297 2179 31331
rect 37289 31297 37323 31331
rect 35817 31229 35851 31263
rect 36737 31229 36771 31263
rect 38117 31093 38151 31127
rect 37381 30753 37415 30787
rect 4169 30685 4203 30719
rect 34989 30685 35023 30719
rect 35817 30685 35851 30719
rect 36277 30685 36311 30719
rect 36461 30617 36495 30651
rect 35081 30277 35115 30311
rect 36737 30277 36771 30311
rect 37381 30277 37415 30311
rect 3985 30209 4019 30243
rect 34897 30209 34931 30243
rect 37289 30209 37323 30243
rect 37933 30209 37967 30243
rect 4169 30141 4203 30175
rect 5549 30141 5583 30175
rect 38025 30141 38059 30175
rect 4353 29801 4387 29835
rect 23397 29665 23431 29699
rect 37197 29665 37231 29699
rect 38117 29665 38151 29699
rect 4445 29597 4479 29631
rect 21097 29597 21131 29631
rect 21557 29597 21591 29631
rect 21741 29529 21775 29563
rect 37933 29529 37967 29563
rect 37473 29257 37507 29291
rect 36737 29121 36771 29155
rect 37381 29121 37415 29155
rect 36645 28917 36679 28951
rect 21005 28713 21039 28747
rect 36461 28577 36495 28611
rect 38117 28577 38151 28611
rect 1869 28509 1903 28543
rect 8953 28509 8987 28543
rect 9873 28509 9907 28543
rect 20913 28509 20947 28543
rect 21741 28509 21775 28543
rect 32321 28509 32355 28543
rect 36277 28509 36311 28543
rect 21557 28441 21591 28475
rect 21925 28373 21959 28407
rect 19533 28101 19567 28135
rect 1777 28033 1811 28067
rect 8493 28033 8527 28067
rect 18797 28033 18831 28067
rect 19901 28033 19935 28067
rect 22753 28033 22787 28067
rect 32321 28033 32355 28067
rect 37657 28033 37691 28067
rect 1961 27965 1995 27999
rect 2237 27965 2271 27999
rect 8677 27965 8711 27999
rect 8953 27965 8987 27999
rect 18613 27965 18647 27999
rect 22569 27965 22603 27999
rect 22661 27965 22695 27999
rect 32505 27965 32539 27999
rect 32873 27965 32907 27999
rect 23121 27829 23155 27863
rect 2145 27625 2179 27659
rect 9045 27625 9079 27659
rect 32597 27625 32631 27659
rect 18613 27557 18647 27591
rect 9781 27489 9815 27523
rect 10241 27489 10275 27523
rect 19533 27489 19567 27523
rect 21005 27489 21039 27523
rect 22017 27489 22051 27523
rect 23305 27489 23339 27523
rect 2237 27421 2271 27455
rect 9137 27421 9171 27455
rect 17601 27421 17635 27455
rect 18337 27421 18371 27455
rect 19257 27421 19291 27455
rect 20821 27421 20855 27455
rect 23029 27421 23063 27455
rect 32689 27421 32723 27455
rect 9965 27353 9999 27387
rect 21833 27353 21867 27387
rect 17693 27285 17727 27319
rect 20637 27285 20671 27319
rect 21465 27285 21499 27319
rect 21925 27285 21959 27319
rect 22661 27285 22695 27319
rect 23121 27285 23155 27319
rect 9965 27081 9999 27115
rect 21833 27081 21867 27115
rect 22201 27081 22235 27115
rect 18613 27013 18647 27047
rect 20085 27013 20119 27047
rect 21005 27013 21039 27047
rect 9873 26945 9907 26979
rect 17417 26945 17451 26979
rect 17877 26945 17911 26979
rect 19349 26945 19383 26979
rect 20729 26945 20763 26979
rect 22293 26945 22327 26979
rect 23213 26945 23247 26979
rect 38025 26945 38059 26979
rect 17233 26877 17267 26911
rect 22385 26877 22419 26911
rect 23397 26877 23431 26911
rect 23029 26741 23063 26775
rect 37933 26741 37967 26775
rect 18245 26401 18279 26435
rect 19717 26401 19751 26435
rect 1685 26333 1719 26367
rect 17509 26333 17543 26367
rect 18613 26333 18647 26367
rect 20545 26333 20579 26367
rect 21281 26333 21315 26367
rect 22109 26333 22143 26367
rect 22293 26333 22327 26367
rect 22569 26333 22603 26367
rect 22753 26333 22787 26367
rect 23397 26333 23431 26367
rect 34713 26333 34747 26367
rect 36277 26333 36311 26367
rect 21097 26265 21131 26299
rect 21465 26265 21499 26299
rect 23213 26265 23247 26299
rect 23581 26265 23615 26299
rect 36461 26265 36495 26299
rect 38117 26265 38151 26299
rect 22845 25993 22879 26027
rect 23213 25993 23247 26027
rect 37381 25993 37415 26027
rect 3433 25925 3467 25959
rect 23673 25925 23707 25959
rect 23857 25925 23891 25959
rect 33517 25925 33551 25959
rect 34253 25925 34287 25959
rect 1593 25857 1627 25891
rect 17141 25857 17175 25891
rect 17601 25857 17635 25891
rect 20545 25857 20579 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22753 25857 22787 25891
rect 33425 25857 33459 25891
rect 36553 25857 36587 25891
rect 37289 25857 37323 25891
rect 37933 25857 37967 25891
rect 1777 25789 1811 25823
rect 17049 25789 17083 25823
rect 17785 25789 17819 25823
rect 18061 25789 18095 25823
rect 20269 25789 20303 25823
rect 22661 25789 22695 25823
rect 34069 25789 34103 25823
rect 35817 25789 35851 25823
rect 21925 25653 21959 25687
rect 24041 25653 24075 25687
rect 38025 25653 38059 25687
rect 2053 25449 2087 25483
rect 20729 25449 20763 25483
rect 25237 25381 25271 25415
rect 20085 25313 20119 25347
rect 21281 25313 21315 25347
rect 21465 25313 21499 25347
rect 22569 25313 22603 25347
rect 25697 25313 25731 25347
rect 27537 25313 27571 25347
rect 37933 25313 37967 25347
rect 2145 25245 2179 25279
rect 18613 25245 18647 25279
rect 20269 25245 20303 25279
rect 20361 25245 20395 25279
rect 22753 25245 22787 25279
rect 23581 25245 23615 25279
rect 23765 25245 23799 25279
rect 25053 25245 25087 25279
rect 38117 25245 38151 25279
rect 18061 25177 18095 25211
rect 21557 25177 21591 25211
rect 25881 25177 25915 25211
rect 36277 25177 36311 25211
rect 21925 25109 21959 25143
rect 22661 25109 22695 25143
rect 23121 25109 23155 25143
rect 23673 25109 23707 25143
rect 24317 24905 24351 24939
rect 25881 24905 25915 24939
rect 22201 24837 22235 24871
rect 18429 24769 18463 24803
rect 19717 24769 19751 24803
rect 20545 24769 20579 24803
rect 21833 24769 21867 24803
rect 21926 24769 21960 24803
rect 22063 24769 22097 24803
rect 22317 24769 22351 24803
rect 23121 24769 23155 24803
rect 23213 24769 23247 24803
rect 23397 24769 23431 24803
rect 23489 24769 23523 24803
rect 23949 24769 23983 24803
rect 24777 24769 24811 24803
rect 24961 24769 24995 24803
rect 25789 24769 25823 24803
rect 37841 24769 37875 24803
rect 19073 24701 19107 24735
rect 24041 24701 24075 24735
rect 24869 24701 24903 24735
rect 22937 24633 22971 24667
rect 22477 24565 22511 24599
rect 23949 24565 23983 24599
rect 17417 24293 17451 24327
rect 22017 24293 22051 24327
rect 24409 24293 24443 24327
rect 21097 24225 21131 24259
rect 21189 24225 21223 24259
rect 23398 24225 23432 24259
rect 23581 24225 23615 24259
rect 25513 24225 25547 24259
rect 27353 24225 27387 24259
rect 1961 24157 1995 24191
rect 17233 24157 17267 24191
rect 18061 24157 18095 24191
rect 20085 24157 20119 24191
rect 20177 24157 20211 24191
rect 20361 24157 20395 24191
rect 20453 24157 20487 24191
rect 21005 24157 21039 24191
rect 21281 24157 21315 24191
rect 22017 24157 22051 24191
rect 22201 24157 22235 24191
rect 22569 24157 22603 24191
rect 22753 24157 22787 24191
rect 23489 24157 23523 24191
rect 23673 24157 23707 24191
rect 24685 24157 24719 24191
rect 37841 24157 37875 24191
rect 18613 24089 18647 24123
rect 24409 24089 24443 24123
rect 25697 24089 25731 24123
rect 19901 24021 19935 24055
rect 21465 24021 21499 24055
rect 23213 24021 23247 24055
rect 24593 24021 24627 24055
rect 21097 23817 21131 23851
rect 25697 23817 25731 23851
rect 3709 23749 3743 23783
rect 18429 23749 18463 23783
rect 1869 23681 1903 23715
rect 19073 23681 19107 23715
rect 19993 23681 20027 23715
rect 21005 23681 21039 23715
rect 22109 23681 22143 23715
rect 22198 23684 22232 23718
rect 22293 23681 22327 23715
rect 22477 23681 22511 23715
rect 23305 23681 23339 23715
rect 25605 23681 25639 23715
rect 37289 23681 37323 23715
rect 2053 23613 2087 23647
rect 19717 23613 19751 23647
rect 23213 23613 23247 23647
rect 21833 23477 21867 23511
rect 23029 23477 23063 23511
rect 37381 23477 37415 23511
rect 2605 23273 2639 23307
rect 23029 23273 23063 23307
rect 21925 23137 21959 23171
rect 22661 23137 22695 23171
rect 37197 23137 37231 23171
rect 37933 23137 37967 23171
rect 38117 23137 38151 23171
rect 1869 23069 1903 23103
rect 2697 23069 2731 23103
rect 19533 23069 19567 23103
rect 20637 23069 20671 23103
rect 21833 23069 21867 23103
rect 23121 23069 23155 23103
rect 28181 23069 28215 23103
rect 19901 23001 19935 23035
rect 20913 23001 20947 23035
rect 1961 22933 1995 22967
rect 22201 22933 22235 22967
rect 28273 22933 28307 22967
rect 20729 22729 20763 22763
rect 28365 22661 28399 22695
rect 19441 22593 19475 22627
rect 20453 22593 20487 22627
rect 21833 22593 21867 22627
rect 22017 22593 22051 22627
rect 22477 22593 22511 22627
rect 22661 22593 22695 22627
rect 28181 22593 28215 22627
rect 37565 22593 37599 22627
rect 19625 22525 19659 22559
rect 30021 22525 30055 22559
rect 22017 22389 22051 22423
rect 22569 22389 22603 22423
rect 36553 22389 36587 22423
rect 37657 22389 37691 22423
rect 22477 22185 22511 22219
rect 22569 22049 22603 22083
rect 36277 22049 36311 22083
rect 38117 22049 38151 22083
rect 19717 21981 19751 22015
rect 20177 21981 20211 22015
rect 22050 21981 22084 22015
rect 19441 21913 19475 21947
rect 36461 21913 36495 21947
rect 21925 21845 21959 21879
rect 22109 21845 22143 21879
rect 19717 21505 19751 21539
rect 22017 21505 22051 21539
rect 23029 21505 23063 21539
rect 37473 21505 37507 21539
rect 21925 21437 21959 21471
rect 22937 21437 22971 21471
rect 22385 21369 22419 21403
rect 23397 21369 23431 21403
rect 19809 21301 19843 21335
rect 36553 21301 36587 21335
rect 37565 21301 37599 21335
rect 19993 20961 20027 20995
rect 22385 20961 22419 20995
rect 36277 20961 36311 20995
rect 36461 20961 36495 20995
rect 38117 20961 38151 20995
rect 22477 20893 22511 20927
rect 24593 20893 24627 20927
rect 20177 20825 20211 20859
rect 21833 20825 21867 20859
rect 22845 20757 22879 20791
rect 24501 20757 24535 20791
rect 23029 20553 23063 20587
rect 23213 20553 23247 20587
rect 23121 20485 23155 20519
rect 23397 20485 23431 20519
rect 24225 20485 24259 20519
rect 2237 20417 2271 20451
rect 2881 20417 2915 20451
rect 22017 20417 22051 20451
rect 24041 20417 24075 20451
rect 37473 20417 37507 20451
rect 25881 20349 25915 20383
rect 22845 20281 22879 20315
rect 1593 20213 1627 20247
rect 2145 20213 2179 20247
rect 2789 20213 2823 20247
rect 22109 20213 22143 20247
rect 37565 20213 37599 20247
rect 1593 19873 1627 19907
rect 1869 19873 1903 19907
rect 22017 19873 22051 19907
rect 22201 19873 22235 19907
rect 24409 19873 24443 19907
rect 37197 19873 37231 19907
rect 37933 19873 37967 19907
rect 1409 19805 1443 19839
rect 21373 19805 21407 19839
rect 31769 19805 31803 19839
rect 38117 19805 38151 19839
rect 23857 19737 23891 19771
rect 24593 19737 24627 19771
rect 26249 19737 26283 19771
rect 21557 19669 21591 19703
rect 31861 19669 31895 19703
rect 24501 19465 24535 19499
rect 1869 19397 1903 19431
rect 32321 19397 32355 19431
rect 1685 19329 1719 19363
rect 22109 19329 22143 19363
rect 23949 19329 23983 19363
rect 24409 19329 24443 19363
rect 37841 19329 37875 19363
rect 2145 19261 2179 19295
rect 22293 19261 22327 19295
rect 31585 19261 31619 19295
rect 32137 19261 32171 19295
rect 32597 19261 32631 19295
rect 1685 18921 1719 18955
rect 21833 18785 21867 18819
rect 20729 18717 20763 18751
rect 21373 18717 21407 18751
rect 20821 18649 20855 18683
rect 21557 18649 21591 18683
rect 22293 18377 22327 18411
rect 22201 18241 22235 18275
rect 26985 18241 27019 18275
rect 1593 18037 1627 18071
rect 27077 18037 27111 18071
rect 27629 18037 27663 18071
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 27077 17697 27111 17731
rect 27261 17697 27295 17731
rect 1593 17561 1627 17595
rect 28917 17561 28951 17595
rect 1961 17289 1995 17323
rect 28365 17221 28399 17255
rect 29101 17221 29135 17255
rect 2053 17153 2087 17187
rect 28273 17153 28307 17187
rect 28917 17085 28951 17119
rect 30757 17085 30791 17119
rect 3617 16949 3651 16983
rect 37841 16949 37875 16983
rect 29561 16745 29595 16779
rect 37657 16609 37691 16643
rect 38117 16609 38151 16643
rect 2145 16541 2179 16575
rect 2789 16541 2823 16575
rect 3801 16541 3835 16575
rect 37933 16473 37967 16507
rect 2053 16405 2087 16439
rect 3893 16405 3927 16439
rect 37565 16201 37599 16235
rect 3249 16133 3283 16167
rect 4077 16133 4111 16167
rect 3433 16065 3467 16099
rect 3893 16065 3927 16099
rect 37473 16065 37507 16099
rect 1593 15997 1627 16031
rect 4353 15997 4387 16031
rect 2789 15521 2823 15555
rect 1409 15453 1443 15487
rect 3985 15453 4019 15487
rect 37841 15453 37875 15487
rect 1593 15317 1627 15351
rect 3893 15317 3927 15351
rect 4261 15045 4295 15079
rect 2053 14977 2087 15011
rect 4445 14977 4479 15011
rect 37473 14977 37507 15011
rect 2881 14909 2915 14943
rect 1961 14773 1995 14807
rect 19809 14773 19843 14807
rect 37565 14773 37599 14807
rect 3065 14433 3099 14467
rect 19809 14433 19843 14467
rect 37197 14433 37231 14467
rect 37933 14433 37967 14467
rect 38117 14433 38151 14467
rect 1409 14365 1443 14399
rect 3249 14365 3283 14399
rect 3801 14365 3835 14399
rect 19993 14297 20027 14331
rect 21649 14297 21683 14331
rect 19441 14025 19475 14059
rect 19349 13889 19383 13923
rect 1869 13821 1903 13855
rect 3525 13821 3559 13855
rect 3709 13821 3743 13855
rect 37841 13685 37875 13719
rect 2605 13481 2639 13515
rect 37197 13345 37231 13379
rect 38117 13345 38151 13379
rect 1593 13277 1627 13311
rect 2697 13277 2731 13311
rect 37933 13209 37967 13243
rect 37565 12937 37599 12971
rect 2053 12801 2087 12835
rect 2697 12801 2731 12835
rect 37473 12801 37507 12835
rect 1961 12597 1995 12631
rect 1409 12257 1443 12291
rect 1593 12257 1627 12291
rect 2789 12257 2823 12291
rect 37197 12257 37231 12291
rect 36277 12189 36311 12223
rect 36461 12121 36495 12155
rect 37565 11713 37599 11747
rect 1685 11645 1719 11679
rect 1869 11645 1903 11679
rect 2789 11645 2823 11679
rect 36553 11509 36587 11543
rect 37657 11509 37691 11543
rect 2053 11305 2087 11339
rect 35817 11305 35851 11339
rect 36277 11169 36311 11203
rect 36461 11169 36495 11203
rect 38117 11169 38151 11203
rect 2145 11101 2179 11135
rect 19717 11101 19751 11135
rect 20269 11033 20303 11067
rect 37565 10761 37599 10795
rect 1685 10625 1719 10659
rect 6561 10625 6595 10659
rect 37473 10625 37507 10659
rect 6469 10421 6503 10455
rect 36553 10421 36587 10455
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 36277 10081 36311 10115
rect 38117 10081 38151 10115
rect 5457 10013 5491 10047
rect 5917 10013 5951 10047
rect 36461 9945 36495 9979
rect 36645 9673 36679 9707
rect 36737 9537 36771 9571
rect 37381 9537 37415 9571
rect 1593 9333 1627 9367
rect 37473 9333 37507 9367
rect 1409 8993 1443 9027
rect 1869 8993 1903 9027
rect 37197 8993 37231 9027
rect 37933 8993 37967 9027
rect 38117 8925 38151 8959
rect 1593 8857 1627 8891
rect 1961 8585 1995 8619
rect 2053 8449 2087 8483
rect 2697 8449 2731 8483
rect 19993 8449 20027 8483
rect 37841 8449 37875 8483
rect 7941 8381 7975 8415
rect 9597 8381 9631 8415
rect 9781 8381 9815 8415
rect 2605 8313 2639 8347
rect 3157 8245 3191 8279
rect 20085 8245 20119 8279
rect 8125 8041 8159 8075
rect 9045 8041 9079 8075
rect 3065 7905 3099 7939
rect 3249 7905 3283 7939
rect 20637 7905 20671 7939
rect 22017 7905 22051 7939
rect 9137 7837 9171 7871
rect 20453 7837 20487 7871
rect 1409 7769 1443 7803
rect 9137 7361 9171 7395
rect 20545 7361 20579 7395
rect 9229 7157 9263 7191
rect 9781 7157 9815 7191
rect 9413 6817 9447 6851
rect 9873 6817 9907 6851
rect 1593 6749 1627 6783
rect 9229 6749 9263 6783
rect 1593 6273 1627 6307
rect 1777 6205 1811 6239
rect 2053 6205 2087 6239
rect 1961 5865 1995 5899
rect 2053 5661 2087 5695
rect 10517 4981 10551 5015
rect 17785 4981 17819 5015
rect 37841 4981 37875 5015
rect 1777 4641 1811 4675
rect 10425 4641 10459 4675
rect 11069 4641 11103 4675
rect 37197 4641 37231 4675
rect 38117 4641 38151 4675
rect 2973 4573 3007 4607
rect 17877 4573 17911 4607
rect 18613 4573 18647 4607
rect 19441 4573 19475 4607
rect 20729 4573 20763 4607
rect 10609 4505 10643 4539
rect 37933 4505 37967 4539
rect 18521 4437 18555 4471
rect 20821 4437 20855 4471
rect 10517 4233 10551 4267
rect 37565 4233 37599 4267
rect 17969 4165 18003 4199
rect 2881 4097 2915 4131
rect 9965 4097 9999 4131
rect 10425 4097 10459 4131
rect 17785 4097 17819 4131
rect 20637 4097 20671 4131
rect 34989 4097 35023 4131
rect 36369 4097 36403 4131
rect 37473 4097 37507 4131
rect 3065 4029 3099 4063
rect 3985 4029 4019 4063
rect 18245 4029 18279 4063
rect 1685 3893 1719 3927
rect 5365 3893 5399 3927
rect 9137 3893 9171 3927
rect 9873 3893 9907 3927
rect 20729 3893 20763 3927
rect 21833 3893 21867 3927
rect 32321 3893 32355 3927
rect 32965 3893 32999 3927
rect 34069 3893 34103 3927
rect 35081 3893 35115 3927
rect 35633 3893 35667 3927
rect 36461 3893 36495 3927
rect 3893 3689 3927 3723
rect 19993 3689 20027 3723
rect 35357 3621 35391 3655
rect 2789 3553 2823 3587
rect 3249 3553 3283 3587
rect 6469 3553 6503 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9597 3553 9631 3587
rect 15669 3553 15703 3587
rect 17969 3553 18003 3587
rect 20821 3553 20855 3587
rect 21281 3553 21315 3587
rect 31585 3553 31619 3587
rect 36829 3553 36863 3587
rect 37841 3553 37875 3587
rect 3985 3485 4019 3519
rect 8125 3485 8159 3519
rect 14381 3485 14415 3519
rect 16129 3485 16163 3519
rect 18429 3485 18463 3519
rect 19257 3485 19291 3519
rect 20177 3485 20211 3519
rect 20637 3485 20671 3519
rect 31033 3485 31067 3519
rect 33333 3485 33367 3519
rect 33977 3485 34011 3519
rect 38025 3485 38059 3519
rect 3065 3417 3099 3451
rect 4629 3417 4663 3451
rect 6285 3417 6319 3451
rect 17785 3417 17819 3451
rect 31217 3417 31251 3451
rect 35173 3417 35207 3451
rect 18521 3349 18555 3383
rect 19349 3349 19383 3383
rect 33425 3349 33459 3383
rect 34069 3349 34103 3383
rect 2697 3145 2731 3179
rect 30849 3145 30883 3179
rect 37749 3145 37783 3179
rect 19165 3077 19199 3111
rect 22017 3077 22051 3111
rect 23673 3077 23707 3111
rect 32781 3077 32815 3111
rect 35081 3077 35115 3111
rect 38025 3077 38059 3111
rect 2145 3009 2179 3043
rect 2605 3009 2639 3043
rect 5641 3009 5675 3043
rect 5733 3009 5767 3043
rect 8677 3009 8711 3043
rect 14289 3009 14323 3043
rect 18981 3009 19015 3043
rect 21833 3009 21867 3043
rect 30757 3009 30791 3043
rect 31401 3009 31435 3043
rect 32597 3009 32631 3043
rect 34897 3009 34931 3043
rect 3341 2941 3375 2975
rect 4997 2941 5031 2975
rect 5181 2941 5215 2975
rect 6377 2941 6411 2975
rect 6561 2941 6595 2975
rect 6837 2941 6871 2975
rect 8861 2941 8895 2975
rect 9137 2941 9171 2975
rect 11529 2941 11563 2975
rect 11713 2941 11747 2975
rect 11989 2941 12023 2975
rect 14473 2941 14507 2975
rect 14841 2941 14875 2975
rect 16681 2941 16715 2975
rect 16865 2941 16899 2975
rect 17141 2941 17175 2975
rect 19441 2941 19475 2975
rect 33517 2941 33551 2975
rect 35449 2941 35483 2975
rect 2053 2805 2087 2839
rect 31493 2805 31527 2839
rect 4721 2601 4755 2635
rect 6377 2601 6411 2635
rect 8033 2601 8067 2635
rect 10517 2601 10551 2635
rect 14473 2601 14507 2635
rect 16129 2601 16163 2635
rect 16773 2601 16807 2635
rect 17417 2601 17451 2635
rect 18613 2601 18647 2635
rect 21833 2601 21867 2635
rect 31033 2601 31067 2635
rect 37473 2601 37507 2635
rect 3985 2533 4019 2567
rect 5549 2533 5583 2567
rect 9965 2533 9999 2567
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 19533 2465 19567 2499
rect 19993 2465 20027 2499
rect 32321 2465 32355 2499
rect 32505 2465 32539 2499
rect 32873 2465 32907 2499
rect 34713 2465 34747 2499
rect 4077 2397 4111 2431
rect 5641 2397 5675 2431
rect 7941 2397 7975 2431
rect 10425 2397 10459 2431
rect 14381 2397 14415 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 19349 2397 19383 2431
rect 18521 2329 18555 2363
rect 34897 2329 34931 2363
rect 36553 2329 36587 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 3418 37408 3424 37460
rect 3476 37448 3482 37460
rect 7466 37448 7472 37460
rect 3476 37420 7472 37448
rect 3476 37408 3482 37420
rect 7466 37408 7472 37420
rect 7524 37408 7530 37460
rect 9953 37451 10011 37457
rect 9953 37417 9965 37451
rect 9999 37448 10011 37451
rect 22462 37448 22468 37460
rect 9999 37420 22468 37448
rect 9999 37417 10011 37420
rect 9953 37411 10011 37417
rect 22462 37408 22468 37420
rect 22520 37408 22526 37460
rect 33505 37451 33563 37457
rect 33505 37417 33517 37451
rect 33551 37448 33563 37451
rect 36170 37448 36176 37460
rect 33551 37420 36176 37448
rect 33551 37417 33563 37420
rect 33505 37411 33563 37417
rect 36170 37408 36176 37420
rect 36228 37408 36234 37460
rect 18693 37383 18751 37389
rect 18693 37349 18705 37383
rect 18739 37380 18751 37383
rect 21818 37380 21824 37392
rect 18739 37352 21824 37380
rect 18739 37349 18751 37352
rect 18693 37343 18751 37349
rect 21818 37340 21824 37352
rect 21876 37340 21882 37392
rect 23382 37340 23388 37392
rect 23440 37380 23446 37392
rect 35342 37380 35348 37392
rect 23440 37352 35348 37380
rect 23440 37340 23446 37352
rect 35342 37340 35348 37352
rect 35400 37340 35406 37392
rect 10689 37315 10747 37321
rect 10689 37281 10701 37315
rect 10735 37312 10747 37315
rect 11422 37312 11428 37324
rect 10735 37284 11428 37312
rect 10735 37281 10747 37284
rect 10689 37275 10747 37281
rect 11422 37272 11428 37284
rect 11480 37272 11486 37324
rect 11698 37272 11704 37324
rect 11756 37312 11762 37324
rect 11977 37315 12035 37321
rect 11977 37312 11989 37315
rect 11756 37284 11989 37312
rect 11756 37272 11762 37284
rect 11977 37281 11989 37284
rect 12023 37281 12035 37315
rect 15194 37312 15200 37324
rect 15155 37284 15200 37312
rect 11977 37275 12035 37281
rect 15194 37272 15200 37284
rect 15252 37272 15258 37324
rect 19978 37312 19984 37324
rect 19939 37284 19984 37312
rect 19978 37272 19984 37284
rect 20036 37272 20042 37324
rect 22005 37315 22063 37321
rect 22005 37281 22017 37315
rect 22051 37312 22063 37315
rect 22554 37312 22560 37324
rect 22051 37284 22560 37312
rect 22051 37281 22063 37284
rect 22005 37275 22063 37281
rect 22554 37272 22560 37284
rect 22612 37272 22618 37324
rect 34149 37315 34207 37321
rect 34149 37281 34161 37315
rect 34195 37312 34207 37315
rect 34790 37312 34796 37324
rect 34195 37284 34796 37312
rect 34195 37281 34207 37284
rect 34149 37275 34207 37281
rect 34790 37272 34796 37284
rect 34848 37272 34854 37324
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 2314 37244 2320 37256
rect 2275 37216 2320 37244
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 3418 37204 3424 37256
rect 3476 37244 3482 37256
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 3476 37216 3801 37244
rect 3476 37204 3482 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 6454 37204 6460 37256
rect 6512 37244 6518 37256
rect 6549 37247 6607 37253
rect 6549 37244 6561 37247
rect 6512 37216 6561 37244
rect 6512 37204 6518 37216
rect 6549 37213 6561 37216
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 7742 37204 7748 37256
rect 7800 37244 7806 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7800 37216 7849 37244
rect 7800 37204 7806 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 11514 37244 11520 37256
rect 11475 37216 11520 37244
rect 9861 37207 9919 37213
rect 11514 37204 11520 37216
rect 11572 37204 11578 37256
rect 14090 37244 14096 37256
rect 14051 37216 14096 37244
rect 14090 37204 14096 37216
rect 14148 37204 14154 37256
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15013 37247 15071 37253
rect 15013 37244 15025 37247
rect 14884 37216 15025 37244
rect 14884 37204 14890 37216
rect 15013 37213 15025 37216
rect 15059 37213 15071 37247
rect 15013 37207 15071 37213
rect 17494 37204 17500 37256
rect 17552 37244 17558 37256
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17552 37216 17601 37244
rect 17552 37204 17558 37216
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 19426 37244 19432 37256
rect 19387 37216 19432 37244
rect 17589 37207 17647 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 20806 37204 20812 37256
rect 20864 37244 20870 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 20864 37216 22753 37244
rect 20864 37204 20870 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 23566 37244 23572 37256
rect 23527 37216 23572 37244
rect 22741 37207 22799 37213
rect 23566 37204 23572 37216
rect 23624 37204 23630 37256
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 7926 37176 7932 37188
rect 1596 37148 7932 37176
rect 1596 37117 1624 37148
rect 7926 37136 7932 37148
rect 7984 37136 7990 37188
rect 8036 37148 10824 37176
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37077 1639 37111
rect 6730 37108 6736 37120
rect 6691 37080 6736 37108
rect 1581 37071 1639 37077
rect 6730 37068 6736 37080
rect 6788 37068 6794 37120
rect 8036 37117 8064 37148
rect 8021 37111 8079 37117
rect 8021 37077 8033 37111
rect 8067 37077 8079 37111
rect 10796 37108 10824 37148
rect 10870 37136 10876 37188
rect 10928 37176 10934 37188
rect 11701 37179 11759 37185
rect 11701 37176 11713 37179
rect 10928 37148 11713 37176
rect 10928 37136 10934 37148
rect 11701 37145 11713 37148
rect 11747 37145 11759 37179
rect 11701 37139 11759 37145
rect 19613 37179 19671 37185
rect 19613 37145 19625 37179
rect 19659 37176 19671 37179
rect 19978 37176 19984 37188
rect 19659 37148 19984 37176
rect 19659 37145 19671 37148
rect 19613 37139 19671 37145
rect 19978 37136 19984 37148
rect 20036 37136 20042 37188
rect 22094 37136 22100 37188
rect 22152 37176 22158 37188
rect 24596 37176 24624 37207
rect 25866 37204 25872 37256
rect 25924 37244 25930 37256
rect 25961 37247 26019 37253
rect 25961 37244 25973 37247
rect 25924 37216 25973 37244
rect 25924 37204 25930 37216
rect 25961 37213 25973 37216
rect 26007 37213 26019 37247
rect 28074 37244 28080 37256
rect 28035 37216 28080 37244
rect 25961 37207 26019 37213
rect 28074 37204 28080 37216
rect 28132 37204 28138 37256
rect 28534 37244 28540 37256
rect 28495 37216 28540 37244
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 33836 37216 34897 37244
rect 33836 37204 33842 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 36722 37244 36728 37256
rect 36683 37216 36728 37244
rect 34885 37207 34943 37213
rect 36722 37204 36728 37216
rect 36780 37204 36786 37256
rect 36814 37204 36820 37256
rect 36872 37244 36878 37256
rect 37369 37247 37427 37253
rect 37369 37244 37381 37247
rect 36872 37216 37381 37244
rect 36872 37204 36878 37216
rect 37369 37213 37381 37216
rect 37415 37213 37427 37247
rect 37369 37207 37427 37213
rect 22152 37148 24624 37176
rect 35069 37179 35127 37185
rect 22152 37136 22158 37148
rect 35069 37145 35081 37179
rect 35115 37176 35127 37179
rect 35342 37176 35348 37188
rect 35115 37148 35348 37176
rect 35115 37145 35127 37148
rect 35069 37139 35127 37145
rect 35342 37136 35348 37148
rect 35400 37136 35406 37188
rect 12342 37108 12348 37120
rect 10796 37080 12348 37108
rect 8021 37071 8079 37077
rect 12342 37068 12348 37080
rect 12400 37068 12406 37120
rect 12434 37068 12440 37120
rect 12492 37108 12498 37120
rect 17402 37108 17408 37120
rect 12492 37080 17408 37108
rect 12492 37068 12498 37080
rect 17402 37068 17408 37080
rect 17460 37068 17466 37120
rect 22833 37111 22891 37117
rect 22833 37077 22845 37111
rect 22879 37108 22891 37111
rect 24302 37108 24308 37120
rect 22879 37080 24308 37108
rect 22879 37077 22891 37080
rect 22833 37071 22891 37077
rect 24302 37068 24308 37080
rect 24360 37068 24366 37120
rect 24394 37068 24400 37120
rect 24452 37108 24458 37120
rect 24452 37080 24497 37108
rect 24452 37068 24458 37080
rect 27890 37068 27896 37120
rect 27948 37108 27954 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27948 37080 27997 37108
rect 27948 37068 27954 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 37458 37108 37464 37120
rect 37419 37080 37464 37108
rect 27985 37071 28043 37077
rect 37458 37068 37464 37080
rect 37516 37068 37522 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 10870 36904 10876 36916
rect 10831 36876 10876 36904
rect 10870 36864 10876 36876
rect 10928 36864 10934 36916
rect 12342 36864 12348 36916
rect 12400 36904 12406 36916
rect 19889 36907 19947 36913
rect 12400 36876 19472 36904
rect 12400 36864 12406 36876
rect 6730 36796 6736 36848
rect 6788 36836 6794 36848
rect 11514 36836 11520 36848
rect 6788 36808 7880 36836
rect 6788 36796 6794 36808
rect 14 36728 20 36780
rect 72 36768 78 36780
rect 1397 36771 1455 36777
rect 1397 36768 1409 36771
rect 72 36740 1409 36768
rect 72 36728 78 36740
rect 1397 36737 1409 36740
rect 1443 36737 1455 36771
rect 1397 36731 1455 36737
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36737 2835 36771
rect 3418 36768 3424 36780
rect 3379 36740 3424 36768
rect 2777 36731 2835 36737
rect 2792 36632 2820 36731
rect 3418 36728 3424 36740
rect 3476 36728 3482 36780
rect 3605 36703 3663 36709
rect 3605 36669 3617 36703
rect 3651 36700 3663 36703
rect 3878 36700 3884 36712
rect 3651 36672 3884 36700
rect 3651 36669 3663 36672
rect 3605 36663 3663 36669
rect 3878 36660 3884 36672
rect 3936 36660 3942 36712
rect 4154 36700 4160 36712
rect 4115 36672 4160 36700
rect 4154 36660 4160 36672
rect 4212 36660 4218 36712
rect 7742 36632 7748 36644
rect 2792 36604 7748 36632
rect 7742 36592 7748 36604
rect 7800 36592 7806 36644
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 1854 36564 1860 36576
rect 1627 36536 1860 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 1854 36524 1860 36536
rect 1912 36524 1918 36576
rect 2685 36567 2743 36573
rect 2685 36533 2697 36567
rect 2731 36564 2743 36567
rect 3050 36564 3056 36576
rect 2731 36536 3056 36564
rect 2731 36533 2743 36536
rect 2685 36527 2743 36533
rect 3050 36524 3056 36536
rect 3108 36524 3114 36576
rect 7852 36564 7880 36808
rect 10336 36808 11520 36836
rect 10336 36777 10364 36808
rect 11514 36796 11520 36808
rect 11572 36796 11578 36848
rect 10321 36771 10379 36777
rect 10321 36737 10333 36771
rect 10367 36737 10379 36771
rect 10778 36768 10784 36780
rect 10739 36740 10784 36768
rect 10321 36731 10379 36737
rect 10778 36728 10784 36740
rect 10836 36728 10842 36780
rect 13633 36771 13691 36777
rect 13633 36737 13645 36771
rect 13679 36768 13691 36771
rect 14090 36768 14096 36780
rect 13679 36740 14096 36768
rect 13679 36737 13691 36740
rect 13633 36731 13691 36737
rect 14090 36728 14096 36740
rect 14148 36728 14154 36780
rect 17494 36768 17500 36780
rect 17455 36740 17500 36768
rect 17494 36728 17500 36740
rect 17552 36728 17558 36780
rect 12250 36700 12256 36712
rect 12211 36672 12256 36700
rect 12250 36660 12256 36672
rect 12308 36660 12314 36712
rect 12618 36660 12624 36712
rect 12676 36700 12682 36712
rect 13449 36703 13507 36709
rect 13449 36700 13461 36703
rect 12676 36672 13461 36700
rect 12676 36660 12682 36672
rect 13449 36669 13461 36672
rect 13495 36669 13507 36703
rect 17678 36700 17684 36712
rect 17639 36672 17684 36700
rect 13449 36663 13507 36669
rect 17678 36660 17684 36672
rect 17736 36660 17742 36712
rect 18046 36700 18052 36712
rect 18007 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 7926 36592 7932 36644
rect 7984 36632 7990 36644
rect 12434 36632 12440 36644
rect 7984 36604 12440 36632
rect 7984 36592 7990 36604
rect 12434 36592 12440 36604
rect 12492 36592 12498 36644
rect 19444 36632 19472 36876
rect 19889 36873 19901 36907
rect 19935 36904 19947 36907
rect 19978 36904 19984 36916
rect 19935 36876 19984 36904
rect 19935 36873 19947 36876
rect 19889 36867 19947 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 21726 36864 21732 36916
rect 21784 36904 21790 36916
rect 24394 36904 24400 36916
rect 21784 36876 24400 36904
rect 21784 36864 21790 36876
rect 24394 36864 24400 36876
rect 24452 36864 24458 36916
rect 20533 36839 20591 36845
rect 20533 36805 20545 36839
rect 20579 36836 20591 36839
rect 22005 36839 22063 36845
rect 22005 36836 22017 36839
rect 20579 36808 22017 36836
rect 20579 36805 20591 36808
rect 20533 36799 20591 36805
rect 22005 36805 22017 36808
rect 22051 36805 22063 36839
rect 24302 36836 24308 36848
rect 24263 36808 24308 36836
rect 22005 36799 22063 36805
rect 24302 36796 24308 36808
rect 24360 36796 24366 36848
rect 27890 36836 27896 36848
rect 27851 36808 27896 36836
rect 27890 36796 27896 36808
rect 27948 36796 27954 36848
rect 35069 36839 35127 36845
rect 35069 36805 35081 36839
rect 35115 36836 35127 36839
rect 37458 36836 37464 36848
rect 35115 36808 37464 36836
rect 35115 36805 35127 36808
rect 35069 36799 35127 36805
rect 37458 36796 37464 36808
rect 37516 36796 37522 36848
rect 19981 36771 20039 36777
rect 19981 36737 19993 36771
rect 20027 36768 20039 36771
rect 20441 36771 20499 36777
rect 20441 36768 20453 36771
rect 20027 36740 20453 36768
rect 20027 36737 20039 36740
rect 19981 36731 20039 36737
rect 20441 36737 20453 36740
rect 20487 36768 20499 36771
rect 20806 36768 20812 36780
rect 20487 36740 20812 36768
rect 20487 36737 20499 36740
rect 20441 36731 20499 36737
rect 20806 36728 20812 36740
rect 20864 36728 20870 36780
rect 21269 36771 21327 36777
rect 21269 36737 21281 36771
rect 21315 36768 21327 36771
rect 21358 36768 21364 36780
rect 21315 36740 21364 36768
rect 21315 36737 21327 36740
rect 21269 36731 21327 36737
rect 21358 36728 21364 36740
rect 21416 36728 21422 36780
rect 21818 36768 21824 36780
rect 21779 36740 21824 36768
rect 21818 36728 21824 36740
rect 21876 36728 21882 36780
rect 23566 36728 23572 36780
rect 23624 36768 23630 36780
rect 24121 36771 24179 36777
rect 24121 36768 24133 36771
rect 23624 36740 24133 36768
rect 23624 36728 23630 36740
rect 24121 36737 24133 36740
rect 24167 36737 24179 36771
rect 33778 36768 33784 36780
rect 33739 36740 33784 36768
rect 24121 36731 24179 36737
rect 33778 36728 33784 36740
rect 33836 36728 33842 36780
rect 34790 36728 34796 36780
rect 34848 36768 34854 36780
rect 34885 36771 34943 36777
rect 34885 36768 34897 36771
rect 34848 36740 34897 36768
rect 34848 36728 34854 36740
rect 34885 36737 34897 36740
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 37182 36768 37188 36780
rect 36771 36740 37188 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 37182 36728 37188 36740
rect 37240 36728 37246 36780
rect 37369 36771 37427 36777
rect 37369 36737 37381 36771
rect 37415 36737 37427 36771
rect 37369 36731 37427 36737
rect 20714 36660 20720 36712
rect 20772 36700 20778 36712
rect 22281 36703 22339 36709
rect 22281 36700 22293 36703
rect 20772 36672 22293 36700
rect 20772 36660 20778 36672
rect 22281 36669 22293 36672
rect 22327 36669 22339 36703
rect 22281 36663 22339 36669
rect 24581 36703 24639 36709
rect 24581 36669 24593 36703
rect 24627 36669 24639 36703
rect 24581 36663 24639 36669
rect 27709 36703 27767 36709
rect 27709 36669 27721 36703
rect 27755 36700 27767 36703
rect 28534 36700 28540 36712
rect 27755 36672 28540 36700
rect 27755 36669 27767 36672
rect 27709 36663 27767 36669
rect 23014 36632 23020 36644
rect 19444 36604 23020 36632
rect 23014 36592 23020 36604
rect 23072 36592 23078 36644
rect 23198 36592 23204 36644
rect 23256 36632 23262 36644
rect 24596 36632 24624 36663
rect 28534 36660 28540 36672
rect 28592 36660 28598 36712
rect 29086 36700 29092 36712
rect 29047 36672 29092 36700
rect 29086 36660 29092 36672
rect 29144 36660 29150 36712
rect 23256 36604 24624 36632
rect 23256 36592 23262 36604
rect 24670 36592 24676 36644
rect 24728 36632 24734 36644
rect 37384 36632 37412 36731
rect 24728 36604 37412 36632
rect 24728 36592 24734 36604
rect 21082 36564 21088 36576
rect 7852 36536 21088 36564
rect 21082 36524 21088 36536
rect 21140 36524 21146 36576
rect 21177 36567 21235 36573
rect 21177 36533 21189 36567
rect 21223 36564 21235 36567
rect 22370 36564 22376 36576
rect 21223 36536 22376 36564
rect 21223 36533 21235 36536
rect 21177 36527 21235 36533
rect 22370 36524 22376 36536
rect 22428 36524 22434 36576
rect 34425 36567 34483 36573
rect 34425 36533 34437 36567
rect 34471 36564 34483 36567
rect 36262 36564 36268 36576
rect 34471 36536 36268 36564
rect 34471 36533 34483 36536
rect 34425 36527 34483 36533
rect 36262 36524 36268 36536
rect 36320 36524 36326 36576
rect 36446 36524 36452 36576
rect 36504 36564 36510 36576
rect 37461 36567 37519 36573
rect 37461 36564 37473 36567
rect 36504 36536 37473 36564
rect 36504 36524 36510 36536
rect 37461 36533 37473 36536
rect 37507 36533 37519 36567
rect 37461 36527 37519 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 3878 36360 3884 36372
rect 3839 36332 3884 36360
rect 3878 36320 3884 36332
rect 3936 36320 3942 36372
rect 7742 36320 7748 36372
rect 7800 36360 7806 36372
rect 10778 36360 10784 36372
rect 7800 36332 10784 36360
rect 7800 36320 7806 36332
rect 10778 36320 10784 36332
rect 10836 36320 10842 36372
rect 12618 36360 12624 36372
rect 12579 36332 12624 36360
rect 12618 36320 12624 36332
rect 12676 36320 12682 36372
rect 17678 36360 17684 36372
rect 17639 36332 17684 36360
rect 17678 36320 17684 36332
rect 17736 36320 17742 36372
rect 19426 36320 19432 36372
rect 19484 36360 19490 36372
rect 19613 36363 19671 36369
rect 19613 36360 19625 36363
rect 19484 36332 19625 36360
rect 19484 36320 19490 36332
rect 19613 36329 19625 36332
rect 19659 36329 19671 36363
rect 19613 36323 19671 36329
rect 21358 36320 21364 36372
rect 21416 36360 21422 36372
rect 24670 36360 24676 36372
rect 21416 36332 24676 36360
rect 21416 36320 21422 36332
rect 24670 36320 24676 36332
rect 24728 36320 24734 36372
rect 35069 36363 35127 36369
rect 35069 36329 35081 36363
rect 35115 36360 35127 36363
rect 35342 36360 35348 36372
rect 35115 36332 35348 36360
rect 35115 36329 35127 36332
rect 35069 36323 35127 36329
rect 35342 36320 35348 36332
rect 35400 36320 35406 36372
rect 2314 36252 2320 36304
rect 2372 36292 2378 36304
rect 2372 36264 3280 36292
rect 2372 36252 2378 36264
rect 1302 36184 1308 36236
rect 1360 36224 1366 36236
rect 1397 36227 1455 36233
rect 1397 36224 1409 36227
rect 1360 36196 1409 36224
rect 1360 36184 1366 36196
rect 1397 36193 1409 36196
rect 1443 36193 1455 36227
rect 3050 36224 3056 36236
rect 3011 36196 3056 36224
rect 1397 36187 1455 36193
rect 3050 36184 3056 36196
rect 3108 36184 3114 36236
rect 3252 36233 3280 36264
rect 21266 36252 21272 36304
rect 21324 36252 21330 36304
rect 36814 36292 36820 36304
rect 25240 36264 36820 36292
rect 3237 36227 3295 36233
rect 3237 36193 3249 36227
rect 3283 36193 3295 36227
rect 3237 36187 3295 36193
rect 7466 36184 7472 36236
rect 7524 36224 7530 36236
rect 10229 36227 10287 36233
rect 10229 36224 10241 36227
rect 7524 36196 10241 36224
rect 7524 36184 7530 36196
rect 10229 36193 10241 36196
rect 10275 36193 10287 36227
rect 10229 36187 10287 36193
rect 11422 36184 11428 36236
rect 11480 36224 11486 36236
rect 12069 36227 12127 36233
rect 12069 36224 12081 36227
rect 11480 36196 12081 36224
rect 11480 36184 11486 36196
rect 12069 36193 12081 36196
rect 12115 36193 12127 36227
rect 12069 36187 12127 36193
rect 21177 36227 21235 36233
rect 21177 36193 21189 36227
rect 21223 36224 21235 36227
rect 21284 36224 21312 36252
rect 22370 36224 22376 36236
rect 21223 36196 21312 36224
rect 22331 36196 22376 36224
rect 21223 36193 21235 36196
rect 21177 36187 21235 36193
rect 22370 36184 22376 36196
rect 22428 36184 22434 36236
rect 22554 36224 22560 36236
rect 22515 36196 22560 36224
rect 22554 36184 22560 36196
rect 22612 36184 22618 36236
rect 25240 36168 25268 36264
rect 36814 36252 36820 36264
rect 36872 36252 36878 36304
rect 25866 36224 25872 36236
rect 25827 36196 25872 36224
rect 25866 36184 25872 36196
rect 25924 36184 25930 36236
rect 26418 36224 26424 36236
rect 26379 36196 26424 36224
rect 26418 36184 26424 36196
rect 26476 36184 26482 36236
rect 36262 36224 36268 36236
rect 36223 36196 36268 36224
rect 36262 36184 36268 36196
rect 36320 36184 36326 36236
rect 36446 36224 36452 36236
rect 36407 36196 36452 36224
rect 36446 36184 36452 36196
rect 36504 36184 36510 36236
rect 38102 36224 38108 36236
rect 38063 36196 38108 36224
rect 38102 36184 38108 36196
rect 38160 36184 38166 36236
rect 3973 36159 4031 36165
rect 3973 36125 3985 36159
rect 4019 36125 4031 36159
rect 12710 36156 12716 36168
rect 12671 36128 12716 36156
rect 3973 36119 4031 36125
rect 3988 36020 4016 36119
rect 12710 36116 12716 36128
rect 12768 36116 12774 36168
rect 17310 36116 17316 36168
rect 17368 36156 17374 36168
rect 17589 36159 17647 36165
rect 17589 36156 17601 36159
rect 17368 36128 17601 36156
rect 17368 36116 17374 36128
rect 17589 36125 17601 36128
rect 17635 36125 17647 36159
rect 17589 36119 17647 36125
rect 23934 36116 23940 36168
rect 23992 36156 23998 36168
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 23992 36128 24409 36156
rect 23992 36116 23998 36128
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 25222 36156 25228 36168
rect 25183 36128 25228 36156
rect 24397 36119 24455 36125
rect 25222 36116 25228 36128
rect 25280 36116 25286 36168
rect 34149 36159 34207 36165
rect 34149 36125 34161 36159
rect 34195 36156 34207 36159
rect 34882 36156 34888 36168
rect 34195 36128 34888 36156
rect 34195 36125 34207 36128
rect 34149 36119 34207 36125
rect 34882 36116 34888 36128
rect 34940 36116 34946 36168
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36156 35035 36159
rect 35434 36156 35440 36168
rect 35023 36128 35440 36156
rect 35023 36125 35035 36128
rect 34977 36119 35035 36125
rect 35434 36116 35440 36128
rect 35492 36116 35498 36168
rect 35618 36156 35624 36168
rect 35579 36128 35624 36156
rect 35618 36116 35624 36128
rect 35676 36116 35682 36168
rect 11882 36088 11888 36100
rect 11843 36060 11888 36088
rect 11882 36048 11888 36060
rect 11940 36048 11946 36100
rect 25317 36091 25375 36097
rect 11992 36060 16574 36088
rect 11992 36020 12020 36060
rect 3988 35992 12020 36020
rect 16546 36020 16574 36060
rect 25317 36057 25329 36091
rect 25363 36088 25375 36091
rect 26053 36091 26111 36097
rect 26053 36088 26065 36091
rect 25363 36060 26065 36088
rect 25363 36057 25375 36060
rect 25317 36051 25375 36057
rect 26053 36057 26065 36060
rect 26099 36057 26111 36091
rect 26053 36051 26111 36057
rect 21358 36020 21364 36032
rect 16546 35992 21364 36020
rect 21358 35980 21364 35992
rect 21416 35980 21422 36032
rect 35713 36023 35771 36029
rect 35713 35989 35725 36023
rect 35759 36020 35771 36023
rect 36446 36020 36452 36032
rect 35759 35992 36452 36020
rect 35759 35989 35771 35992
rect 35713 35983 35771 35989
rect 36446 35980 36452 35992
rect 36504 35980 36510 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 11609 35819 11667 35825
rect 11609 35785 11621 35819
rect 11655 35816 11667 35819
rect 11882 35816 11888 35828
rect 11655 35788 11888 35816
rect 11655 35785 11667 35788
rect 11609 35779 11667 35785
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 28350 35776 28356 35828
rect 28408 35816 28414 35828
rect 29086 35816 29092 35828
rect 28408 35788 29092 35816
rect 28408 35776 28414 35788
rect 29086 35776 29092 35788
rect 29144 35776 29150 35828
rect 36722 35748 36728 35760
rect 36683 35720 36728 35748
rect 36722 35708 36728 35720
rect 36780 35708 36786 35760
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35680 11759 35683
rect 12710 35680 12716 35692
rect 11747 35652 12716 35680
rect 11747 35649 11759 35652
rect 11701 35643 11759 35649
rect 12710 35640 12716 35652
rect 12768 35640 12774 35692
rect 23934 35680 23940 35692
rect 23895 35652 23940 35680
rect 23934 35640 23940 35652
rect 23992 35640 23998 35692
rect 34882 35680 34888 35692
rect 34843 35652 34888 35680
rect 34882 35640 34888 35652
rect 34940 35640 34946 35692
rect 38010 35680 38016 35692
rect 37971 35652 38016 35680
rect 38010 35640 38016 35652
rect 38068 35640 38074 35692
rect 24121 35615 24179 35621
rect 24121 35581 24133 35615
rect 24167 35612 24179 35615
rect 24486 35612 24492 35624
rect 24167 35584 24492 35612
rect 24167 35581 24179 35584
rect 24121 35575 24179 35581
rect 24486 35572 24492 35584
rect 24544 35572 24550 35624
rect 24578 35572 24584 35624
rect 24636 35612 24642 35624
rect 35069 35615 35127 35621
rect 24636 35584 24681 35612
rect 24636 35572 24642 35584
rect 35069 35581 35081 35615
rect 35115 35612 35127 35615
rect 35526 35612 35532 35624
rect 35115 35584 35532 35612
rect 35115 35581 35127 35584
rect 35069 35575 35127 35581
rect 35526 35572 35532 35584
rect 35584 35572 35590 35624
rect 23290 35436 23296 35488
rect 23348 35476 23354 35488
rect 37921 35479 37979 35485
rect 37921 35476 37933 35479
rect 23348 35448 37933 35476
rect 23348 35436 23354 35448
rect 37921 35445 37933 35448
rect 37967 35445 37979 35479
rect 37921 35439 37979 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 24486 35272 24492 35284
rect 24447 35244 24492 35272
rect 24486 35232 24492 35244
rect 24544 35232 24550 35284
rect 35526 35232 35532 35284
rect 35584 35272 35590 35284
rect 35621 35275 35679 35281
rect 35621 35272 35633 35275
rect 35584 35244 35633 35272
rect 35584 35232 35590 35244
rect 35621 35241 35633 35244
rect 35667 35241 35679 35275
rect 35621 35235 35679 35241
rect 36170 35096 36176 35148
rect 36228 35136 36234 35148
rect 36265 35139 36323 35145
rect 36265 35136 36277 35139
rect 36228 35108 36277 35136
rect 36228 35096 36234 35108
rect 36265 35105 36277 35108
rect 36311 35105 36323 35139
rect 36446 35136 36452 35148
rect 36407 35108 36452 35136
rect 36265 35099 36323 35105
rect 36446 35096 36452 35108
rect 36504 35096 36510 35148
rect 38102 35136 38108 35148
rect 38063 35108 38108 35136
rect 38102 35096 38108 35108
rect 38160 35096 38166 35148
rect 1578 35028 1584 35080
rect 1636 35068 1642 35080
rect 1673 35071 1731 35077
rect 1673 35068 1685 35071
rect 1636 35040 1685 35068
rect 1636 35028 1642 35040
rect 1673 35037 1685 35040
rect 1719 35037 1731 35071
rect 1673 35031 1731 35037
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35068 24639 35071
rect 24670 35068 24676 35080
rect 24627 35040 24676 35068
rect 24627 35037 24639 35040
rect 24581 35031 24639 35037
rect 24670 35028 24676 35040
rect 24728 35068 24734 35080
rect 24728 35040 26234 35068
rect 24728 35028 24734 35040
rect 26206 34932 26234 35040
rect 35434 35028 35440 35080
rect 35492 35068 35498 35080
rect 35529 35071 35587 35077
rect 35529 35068 35541 35071
rect 35492 35040 35541 35068
rect 35492 35028 35498 35040
rect 35529 35037 35541 35040
rect 35575 35037 35587 35071
rect 35529 35031 35587 35037
rect 37458 34932 37464 34944
rect 26206 34904 37464 34932
rect 37458 34892 37464 34904
rect 37516 34892 37522 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 29270 34620 29276 34672
rect 29328 34660 29334 34672
rect 32214 34660 32220 34672
rect 29328 34632 32220 34660
rect 29328 34620 29334 34632
rect 32214 34620 32220 34632
rect 32272 34620 32278 34672
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 27338 34552 27344 34604
rect 27396 34592 27402 34604
rect 29638 34592 29644 34604
rect 27396 34564 29644 34592
rect 27396 34552 27402 34564
rect 29638 34552 29644 34564
rect 29696 34552 29702 34604
rect 37458 34592 37464 34604
rect 37419 34564 37464 34592
rect 37458 34552 37464 34564
rect 37516 34552 37522 34604
rect 1762 34524 1768 34536
rect 1723 34496 1768 34524
rect 1762 34484 1768 34496
rect 1820 34484 1826 34536
rect 2774 34524 2780 34536
rect 2735 34496 2780 34524
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 4614 34484 4620 34536
rect 4672 34524 4678 34536
rect 5534 34524 5540 34536
rect 4672 34496 5540 34524
rect 4672 34484 4678 34496
rect 5534 34484 5540 34496
rect 5592 34484 5598 34536
rect 28258 34484 28264 34536
rect 28316 34524 28322 34536
rect 30926 34524 30932 34536
rect 28316 34496 30932 34524
rect 28316 34484 28322 34496
rect 30926 34484 30932 34496
rect 30984 34484 30990 34536
rect 36446 34484 36452 34536
rect 36504 34524 36510 34536
rect 37553 34527 37611 34533
rect 37553 34524 37565 34527
rect 36504 34496 37565 34524
rect 36504 34484 36510 34496
rect 37553 34493 37565 34496
rect 37599 34493 37611 34527
rect 37553 34487 37611 34493
rect 36262 34348 36268 34400
rect 36320 34388 36326 34400
rect 36541 34391 36599 34397
rect 36541 34388 36553 34391
rect 36320 34360 36553 34388
rect 36320 34348 36326 34360
rect 36541 34357 36553 34360
rect 36587 34357 36599 34391
rect 36541 34351 36599 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1762 34144 1768 34196
rect 1820 34184 1826 34196
rect 2041 34187 2099 34193
rect 2041 34184 2053 34187
rect 1820 34156 2053 34184
rect 1820 34144 1826 34156
rect 2041 34153 2053 34156
rect 2087 34153 2099 34187
rect 2041 34147 2099 34153
rect 36262 34048 36268 34060
rect 36223 34020 36268 34048
rect 36262 34008 36268 34020
rect 36320 34008 36326 34060
rect 36446 34048 36452 34060
rect 36407 34020 36452 34048
rect 36446 34008 36452 34020
rect 36504 34008 36510 34060
rect 38102 34048 38108 34060
rect 38063 34020 38108 34048
rect 38102 34008 38108 34020
rect 38160 34008 38166 34060
rect 2133 33983 2191 33989
rect 2133 33949 2145 33983
rect 2179 33980 2191 33983
rect 17310 33980 17316 33992
rect 2179 33952 17316 33980
rect 2179 33949 2191 33952
rect 2133 33943 2191 33949
rect 17310 33940 17316 33952
rect 17368 33940 17374 33992
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 26421 33575 26479 33581
rect 26421 33541 26433 33575
rect 26467 33572 26479 33575
rect 29270 33572 29276 33584
rect 26467 33544 29276 33572
rect 26467 33541 26479 33544
rect 26421 33535 26479 33541
rect 29270 33532 29276 33544
rect 29328 33532 29334 33584
rect 38010 33504 38016 33516
rect 37971 33476 38016 33504
rect 38010 33464 38016 33476
rect 38068 33464 38074 33516
rect 24578 33436 24584 33448
rect 24539 33408 24584 33436
rect 24578 33396 24584 33408
rect 24636 33396 24642 33448
rect 24762 33436 24768 33448
rect 24723 33408 24768 33436
rect 24762 33396 24768 33408
rect 24820 33396 24826 33448
rect 37826 33368 37832 33380
rect 37787 33340 37832 33368
rect 37826 33328 37832 33340
rect 37884 33328 37890 33380
rect 18598 33300 18604 33312
rect 18559 33272 18604 33300
rect 18598 33260 18604 33272
rect 18656 33260 18662 33312
rect 36538 33300 36544 33312
rect 36499 33272 36544 33300
rect 36538 33260 36544 33272
rect 36596 33260 36602 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 24578 33056 24584 33108
rect 24636 33096 24642 33108
rect 24673 33099 24731 33105
rect 24673 33096 24685 33099
rect 24636 33068 24685 33096
rect 24636 33056 24642 33068
rect 24673 33065 24685 33068
rect 24719 33065 24731 33099
rect 24673 33059 24731 33065
rect 6886 33000 19748 33028
rect 3418 32784 3424 32836
rect 3476 32824 3482 32836
rect 6886 32824 6914 33000
rect 18598 32920 18604 32972
rect 18656 32960 18662 32972
rect 19720 32969 19748 33000
rect 19245 32963 19303 32969
rect 19245 32960 19257 32963
rect 18656 32932 19257 32960
rect 18656 32920 18662 32932
rect 19245 32929 19257 32932
rect 19291 32929 19303 32963
rect 19245 32923 19303 32929
rect 19705 32963 19763 32969
rect 19705 32929 19717 32963
rect 19751 32929 19763 32963
rect 19705 32923 19763 32929
rect 36265 32963 36323 32969
rect 36265 32929 36277 32963
rect 36311 32960 36323 32963
rect 36538 32960 36544 32972
rect 36311 32932 36544 32960
rect 36311 32929 36323 32932
rect 36265 32923 36323 32929
rect 36538 32920 36544 32932
rect 36596 32920 36602 32972
rect 3476 32796 6914 32824
rect 3476 32784 3482 32796
rect 19150 32784 19156 32836
rect 19208 32824 19214 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 19208 32796 19441 32824
rect 19208 32784 19214 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 19429 32787 19487 32793
rect 36449 32827 36507 32833
rect 36449 32793 36461 32827
rect 36495 32824 36507 32827
rect 36630 32824 36636 32836
rect 36495 32796 36636 32824
rect 36495 32793 36507 32796
rect 36449 32787 36507 32793
rect 36630 32784 36636 32796
rect 36688 32784 36694 32836
rect 38102 32824 38108 32836
rect 38063 32796 38108 32824
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 19150 32552 19156 32564
rect 19111 32524 19156 32552
rect 19150 32512 19156 32524
rect 19208 32512 19214 32564
rect 24305 32555 24363 32561
rect 24305 32521 24317 32555
rect 24351 32552 24363 32555
rect 24762 32552 24768 32564
rect 24351 32524 24768 32552
rect 24351 32521 24363 32524
rect 24305 32515 24363 32521
rect 24762 32512 24768 32524
rect 24820 32512 24826 32564
rect 36630 32552 36636 32564
rect 36591 32524 36636 32552
rect 36630 32512 36636 32524
rect 36688 32512 36694 32564
rect 19245 32419 19303 32425
rect 19245 32385 19257 32419
rect 19291 32416 19303 32419
rect 20254 32416 20260 32428
rect 19291 32388 20260 32416
rect 19291 32385 19303 32388
rect 19245 32379 19303 32385
rect 20254 32376 20260 32388
rect 20312 32376 20318 32428
rect 21266 32376 21272 32428
rect 21324 32416 21330 32428
rect 24213 32419 24271 32425
rect 24213 32416 24225 32419
rect 21324 32388 24225 32416
rect 21324 32376 21330 32388
rect 24213 32385 24225 32388
rect 24259 32385 24271 32419
rect 36725 32419 36783 32425
rect 36725 32416 36737 32419
rect 24213 32379 24271 32385
rect 26206 32388 36737 32416
rect 12710 32308 12716 32360
rect 12768 32348 12774 32360
rect 17218 32348 17224 32360
rect 12768 32320 17224 32348
rect 12768 32308 12774 32320
rect 17218 32308 17224 32320
rect 17276 32348 17282 32360
rect 26206 32348 26234 32388
rect 36725 32385 36737 32388
rect 36771 32385 36783 32419
rect 36725 32379 36783 32385
rect 37369 32419 37427 32425
rect 37369 32385 37381 32419
rect 37415 32416 37427 32419
rect 37642 32416 37648 32428
rect 37415 32388 37648 32416
rect 37415 32385 37427 32388
rect 37369 32379 37427 32385
rect 17276 32320 26234 32348
rect 36740 32348 36768 32379
rect 37642 32376 37648 32388
rect 37700 32376 37706 32428
rect 37918 32348 37924 32360
rect 36740 32320 37924 32348
rect 17276 32308 17282 32320
rect 37918 32308 37924 32320
rect 37976 32308 37982 32360
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1673 32215 1731 32221
rect 1673 32212 1685 32215
rect 1452 32184 1685 32212
rect 1452 32172 1458 32184
rect 1673 32181 1685 32184
rect 1719 32181 1731 32215
rect 1673 32175 1731 32181
rect 36081 32215 36139 32221
rect 36081 32181 36093 32215
rect 36127 32212 36139 32215
rect 36262 32212 36268 32224
rect 36127 32184 36268 32212
rect 36127 32181 36139 32184
rect 36081 32175 36139 32181
rect 36262 32172 36268 32184
rect 36320 32172 36326 32224
rect 36446 32172 36452 32224
rect 36504 32212 36510 32224
rect 37461 32215 37519 32221
rect 37461 32212 37473 32215
rect 36504 32184 37473 32212
rect 36504 32172 36510 32184
rect 37461 32181 37473 32184
rect 37507 32181 37519 32215
rect 37461 32175 37519 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 36262 31872 36268 31884
rect 36223 31844 36268 31872
rect 36262 31832 36268 31844
rect 36320 31832 36326 31884
rect 36446 31872 36452 31884
rect 36407 31844 36452 31872
rect 36446 31832 36452 31844
rect 36504 31832 36510 31884
rect 38102 31872 38108 31884
rect 38063 31844 38108 31872
rect 38102 31832 38108 31844
rect 38160 31832 38166 31884
rect 35805 31807 35863 31813
rect 35805 31773 35817 31807
rect 35851 31804 35863 31807
rect 36170 31804 36176 31816
rect 35851 31776 36176 31804
rect 35851 31773 35863 31776
rect 35805 31767 35863 31773
rect 36170 31764 36176 31776
rect 36228 31764 36234 31816
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2041 31467 2099 31473
rect 2041 31464 2053 31467
rect 1636 31436 2053 31464
rect 1636 31424 1642 31436
rect 2041 31433 2053 31436
rect 2087 31433 2099 31467
rect 2041 31427 2099 31433
rect 36541 31399 36599 31405
rect 36541 31365 36553 31399
rect 36587 31396 36599 31399
rect 37369 31399 37427 31405
rect 37369 31396 37381 31399
rect 36587 31368 37381 31396
rect 36587 31365 36599 31368
rect 36541 31359 36599 31365
rect 37369 31365 37381 31368
rect 37415 31365 37427 31399
rect 37369 31359 37427 31365
rect 2130 31328 2136 31340
rect 2091 31300 2136 31328
rect 2130 31288 2136 31300
rect 2188 31288 2194 31340
rect 37277 31331 37335 31337
rect 37277 31297 37289 31331
rect 37323 31328 37335 31331
rect 37458 31328 37464 31340
rect 37323 31300 37464 31328
rect 37323 31297 37335 31300
rect 37277 31291 37335 31297
rect 37458 31288 37464 31300
rect 37516 31288 37522 31340
rect 35802 31260 35808 31272
rect 35763 31232 35808 31260
rect 35802 31220 35808 31232
rect 35860 31220 35866 31272
rect 36170 31220 36176 31272
rect 36228 31260 36234 31272
rect 36725 31263 36783 31269
rect 36725 31260 36737 31263
rect 36228 31232 36737 31260
rect 36228 31220 36234 31232
rect 36725 31229 36737 31232
rect 36771 31229 36783 31263
rect 36725 31223 36783 31229
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 10962 31124 10968 31136
rect 9732 31096 10968 31124
rect 9732 31084 9738 31096
rect 10962 31084 10968 31096
rect 11020 31084 11026 31136
rect 38102 31124 38108 31136
rect 38063 31096 38108 31124
rect 38102 31084 38108 31096
rect 38160 31084 38166 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 37366 30784 37372 30796
rect 37327 30756 37372 30784
rect 37366 30744 37372 30756
rect 37424 30744 37430 30796
rect 4154 30716 4160 30728
rect 4115 30688 4160 30716
rect 4154 30676 4160 30688
rect 4212 30676 4218 30728
rect 34882 30676 34888 30728
rect 34940 30716 34946 30728
rect 34977 30719 35035 30725
rect 34977 30716 34989 30719
rect 34940 30688 34989 30716
rect 34940 30676 34946 30688
rect 34977 30685 34989 30688
rect 35023 30685 35035 30719
rect 34977 30679 35035 30685
rect 35805 30719 35863 30725
rect 35805 30685 35817 30719
rect 35851 30716 35863 30719
rect 36265 30719 36323 30725
rect 36265 30716 36277 30719
rect 35851 30688 36277 30716
rect 35851 30685 35863 30688
rect 35805 30679 35863 30685
rect 36265 30685 36277 30688
rect 36311 30685 36323 30719
rect 36265 30679 36323 30685
rect 36449 30651 36507 30657
rect 36449 30617 36461 30651
rect 36495 30648 36507 30651
rect 37366 30648 37372 30660
rect 36495 30620 37372 30648
rect 36495 30617 36507 30620
rect 36449 30611 36507 30617
rect 37366 30608 37372 30620
rect 37424 30608 37430 30660
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4154 30308 4160 30320
rect 3988 30280 4160 30308
rect 3988 30249 4016 30280
rect 4154 30268 4160 30280
rect 4212 30268 4218 30320
rect 35069 30311 35127 30317
rect 35069 30277 35081 30311
rect 35115 30308 35127 30311
rect 36722 30308 36728 30320
rect 35115 30280 36584 30308
rect 36683 30280 36728 30308
rect 35115 30277 35127 30280
rect 35069 30271 35127 30277
rect 3973 30243 4031 30249
rect 3973 30209 3985 30243
rect 4019 30209 4031 30243
rect 34882 30240 34888 30252
rect 34843 30212 34888 30240
rect 3973 30203 4031 30209
rect 34882 30200 34888 30212
rect 34940 30200 34946 30252
rect 4157 30175 4215 30181
rect 4157 30141 4169 30175
rect 4203 30172 4215 30175
rect 4614 30172 4620 30184
rect 4203 30144 4620 30172
rect 4203 30141 4215 30144
rect 4157 30135 4215 30141
rect 4614 30132 4620 30144
rect 4672 30132 4678 30184
rect 5534 30172 5540 30184
rect 5495 30144 5540 30172
rect 5534 30132 5540 30144
rect 5592 30132 5598 30184
rect 36556 30172 36584 30280
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 37366 30308 37372 30320
rect 37327 30280 37372 30308
rect 37366 30268 37372 30280
rect 37424 30268 37430 30320
rect 37274 30240 37280 30252
rect 37235 30212 37280 30240
rect 37274 30200 37280 30212
rect 37332 30200 37338 30252
rect 37918 30240 37924 30252
rect 37879 30212 37924 30240
rect 37918 30200 37924 30212
rect 37976 30200 37982 30252
rect 38013 30175 38071 30181
rect 38013 30172 38025 30175
rect 36556 30144 38025 30172
rect 38013 30141 38025 30144
rect 38059 30141 38071 30175
rect 38013 30135 38071 30141
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 4341 29835 4399 29841
rect 4341 29801 4353 29835
rect 4387 29832 4399 29835
rect 4614 29832 4620 29844
rect 4387 29804 4620 29832
rect 4387 29801 4399 29804
rect 4341 29795 4399 29801
rect 4614 29792 4620 29804
rect 4672 29792 4678 29844
rect 23382 29696 23388 29708
rect 23343 29668 23388 29696
rect 23382 29656 23388 29668
rect 23440 29656 23446 29708
rect 37182 29696 37188 29708
rect 37143 29668 37188 29696
rect 37182 29656 37188 29668
rect 37240 29656 37246 29708
rect 38102 29696 38108 29708
rect 38063 29668 38108 29696
rect 38102 29656 38108 29668
rect 38160 29656 38166 29708
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29628 4491 29631
rect 4798 29628 4804 29640
rect 4479 29600 4804 29628
rect 4479 29597 4491 29600
rect 4433 29591 4491 29597
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29628 21143 29631
rect 21545 29631 21603 29637
rect 21545 29628 21557 29631
rect 21131 29600 21557 29628
rect 21131 29597 21143 29600
rect 21085 29591 21143 29597
rect 21545 29597 21557 29600
rect 21591 29597 21603 29631
rect 21545 29591 21603 29597
rect 21726 29560 21732 29572
rect 21687 29532 21732 29560
rect 21726 29520 21732 29532
rect 21784 29520 21790 29572
rect 37458 29520 37464 29572
rect 37516 29560 37522 29572
rect 37921 29563 37979 29569
rect 37921 29560 37933 29563
rect 37516 29532 37933 29560
rect 37516 29520 37522 29532
rect 37921 29529 37933 29532
rect 37967 29529 37979 29563
rect 37921 29523 37979 29529
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 37458 29288 37464 29300
rect 37419 29260 37464 29288
rect 37458 29248 37464 29260
rect 37516 29248 37522 29300
rect 36725 29155 36783 29161
rect 36725 29121 36737 29155
rect 36771 29121 36783 29155
rect 36725 29115 36783 29121
rect 36740 29084 36768 29115
rect 37274 29112 37280 29164
rect 37332 29152 37338 29164
rect 37369 29155 37427 29161
rect 37369 29152 37381 29155
rect 37332 29124 37381 29152
rect 37332 29112 37338 29124
rect 37369 29121 37381 29124
rect 37415 29152 37427 29155
rect 37458 29152 37464 29164
rect 37415 29124 37464 29152
rect 37415 29121 37427 29124
rect 37369 29115 37427 29121
rect 37458 29112 37464 29124
rect 37516 29112 37522 29164
rect 37550 29084 37556 29096
rect 36740 29056 37556 29084
rect 37550 29044 37556 29056
rect 37608 29044 37614 29096
rect 36446 28908 36452 28960
rect 36504 28948 36510 28960
rect 36633 28951 36691 28957
rect 36633 28948 36645 28951
rect 36504 28920 36645 28948
rect 36504 28908 36510 28920
rect 36633 28917 36645 28920
rect 36679 28917 36691 28951
rect 36633 28911 36691 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 20993 28747 21051 28753
rect 20993 28713 21005 28747
rect 21039 28744 21051 28747
rect 21726 28744 21732 28756
rect 21039 28716 21732 28744
rect 21039 28713 21051 28716
rect 20993 28707 21051 28713
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 36446 28608 36452 28620
rect 36407 28580 36452 28608
rect 36446 28568 36452 28580
rect 36504 28568 36510 28620
rect 38102 28608 38108 28620
rect 38063 28580 38108 28608
rect 38102 28568 38108 28580
rect 38160 28568 38166 28620
rect 1762 28500 1768 28552
rect 1820 28540 1826 28552
rect 1857 28543 1915 28549
rect 1857 28540 1869 28543
rect 1820 28512 1869 28540
rect 1820 28500 1826 28512
rect 1857 28509 1869 28512
rect 1903 28509 1915 28543
rect 1857 28503 1915 28509
rect 8478 28500 8484 28552
rect 8536 28540 8542 28552
rect 8941 28543 8999 28549
rect 8941 28540 8953 28543
rect 8536 28512 8953 28540
rect 8536 28500 8542 28512
rect 8941 28509 8953 28512
rect 8987 28509 8999 28543
rect 8941 28503 8999 28509
rect 9766 28500 9772 28552
rect 9824 28540 9830 28552
rect 9861 28543 9919 28549
rect 9861 28540 9873 28543
rect 9824 28512 9873 28540
rect 9824 28500 9830 28512
rect 9861 28509 9873 28512
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 18598 28500 18604 28552
rect 18656 28540 18662 28552
rect 20901 28543 20959 28549
rect 20901 28540 20913 28543
rect 18656 28512 20913 28540
rect 18656 28500 18662 28512
rect 20901 28509 20913 28512
rect 20947 28509 20959 28543
rect 20901 28503 20959 28509
rect 21729 28543 21787 28549
rect 21729 28509 21741 28543
rect 21775 28540 21787 28543
rect 21818 28540 21824 28552
rect 21775 28512 21824 28540
rect 21775 28509 21787 28512
rect 21729 28503 21787 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 32306 28540 32312 28552
rect 32267 28512 32312 28540
rect 32306 28500 32312 28512
rect 32364 28500 32370 28552
rect 36262 28540 36268 28552
rect 36223 28512 36268 28540
rect 36262 28500 36268 28512
rect 36320 28500 36326 28552
rect 21542 28472 21548 28484
rect 21503 28444 21548 28472
rect 21542 28432 21548 28444
rect 21600 28432 21606 28484
rect 21910 28404 21916 28416
rect 21871 28376 21916 28404
rect 21910 28364 21916 28376
rect 21968 28364 21974 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 33318 28200 33324 28212
rect 19536 28172 33324 28200
rect 19426 28092 19432 28144
rect 19484 28132 19490 28144
rect 19536 28141 19564 28172
rect 33318 28160 33324 28172
rect 33376 28160 33382 28212
rect 19521 28135 19579 28141
rect 19521 28132 19533 28135
rect 19484 28104 19533 28132
rect 19484 28092 19490 28104
rect 19521 28101 19533 28104
rect 19567 28101 19579 28135
rect 19521 28095 19579 28101
rect 22066 28104 31754 28132
rect 1762 28064 1768 28076
rect 1723 28036 1768 28064
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 8478 28064 8484 28076
rect 8439 28036 8484 28064
rect 8478 28024 8484 28036
rect 8536 28024 8542 28076
rect 18782 28064 18788 28076
rect 18743 28036 18788 28064
rect 18782 28024 18788 28036
rect 18840 28024 18846 28076
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19392 28036 19901 28064
rect 19392 28024 19398 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 22066 28064 22094 28104
rect 31726 28076 31754 28104
rect 19889 28027 19947 28033
rect 21100 28036 22094 28064
rect 1946 27996 1952 28008
rect 1907 27968 1952 27996
rect 1946 27956 1952 27968
rect 2004 27956 2010 28008
rect 2225 27999 2283 28005
rect 2225 27965 2237 27999
rect 2271 27965 2283 27999
rect 8662 27996 8668 28008
rect 8623 27968 8668 27996
rect 2225 27959 2283 27965
rect 1486 27888 1492 27940
rect 1544 27928 1550 27940
rect 2240 27928 2268 27959
rect 8662 27956 8668 27968
rect 8720 27956 8726 28008
rect 8941 27999 8999 28005
rect 8941 27965 8953 27999
rect 8987 27965 8999 27999
rect 8941 27959 8999 27965
rect 1544 27900 2268 27928
rect 1544 27888 1550 27900
rect 8294 27888 8300 27940
rect 8352 27928 8358 27940
rect 8956 27928 8984 27959
rect 18414 27956 18420 28008
rect 18472 27996 18478 28008
rect 18601 27999 18659 28005
rect 18601 27996 18613 27999
rect 18472 27968 18613 27996
rect 18472 27956 18478 27968
rect 18601 27965 18613 27968
rect 18647 27996 18659 27999
rect 21100 27996 21128 28036
rect 22462 28024 22468 28076
rect 22520 28064 22526 28076
rect 22741 28067 22799 28073
rect 22741 28064 22753 28067
rect 22520 28036 22753 28064
rect 22520 28024 22526 28036
rect 22741 28033 22753 28036
rect 22787 28033 22799 28067
rect 31726 28036 31760 28076
rect 22741 28027 22799 28033
rect 31754 28024 31760 28036
rect 31812 28024 31818 28076
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 36262 28024 36268 28076
rect 36320 28064 36326 28076
rect 37645 28067 37703 28073
rect 37645 28064 37657 28067
rect 36320 28036 37657 28064
rect 36320 28024 36326 28036
rect 37645 28033 37657 28036
rect 37691 28033 37703 28067
rect 37645 28027 37703 28033
rect 18647 27968 21128 27996
rect 22557 27999 22615 28005
rect 18647 27965 18659 27968
rect 18601 27959 18659 27965
rect 22557 27965 22569 27999
rect 22603 27965 22615 27999
rect 22557 27959 22615 27965
rect 8352 27900 8984 27928
rect 22572 27928 22600 27959
rect 22646 27956 22652 28008
rect 22704 27996 22710 28008
rect 32490 27996 32496 28008
rect 22704 27968 22749 27996
rect 32451 27968 32496 27996
rect 22704 27956 22710 27968
rect 32490 27956 32496 27968
rect 32548 27956 32554 28008
rect 32858 27996 32864 28008
rect 32819 27968 32864 27996
rect 32858 27956 32864 27968
rect 32916 27956 32922 28008
rect 23290 27928 23296 27940
rect 22572 27900 23296 27928
rect 8352 27888 8358 27900
rect 23290 27888 23296 27900
rect 23348 27888 23354 27940
rect 23109 27863 23167 27869
rect 23109 27829 23121 27863
rect 23155 27860 23167 27863
rect 23198 27860 23204 27872
rect 23155 27832 23204 27860
rect 23155 27829 23167 27832
rect 23109 27823 23167 27829
rect 23198 27820 23204 27832
rect 23256 27820 23262 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1946 27616 1952 27668
rect 2004 27656 2010 27668
rect 2133 27659 2191 27665
rect 2133 27656 2145 27659
rect 2004 27628 2145 27656
rect 2004 27616 2010 27628
rect 2133 27625 2145 27628
rect 2179 27625 2191 27659
rect 2133 27619 2191 27625
rect 8662 27616 8668 27668
rect 8720 27656 8726 27668
rect 9033 27659 9091 27665
rect 9033 27656 9045 27659
rect 8720 27628 9045 27656
rect 8720 27616 8726 27628
rect 9033 27625 9045 27628
rect 9079 27625 9091 27659
rect 9033 27619 9091 27625
rect 32490 27616 32496 27668
rect 32548 27656 32554 27668
rect 32585 27659 32643 27665
rect 32585 27656 32597 27659
rect 32548 27628 32597 27656
rect 32548 27616 32554 27628
rect 32585 27625 32597 27628
rect 32631 27625 32643 27659
rect 32585 27619 32643 27625
rect 18598 27588 18604 27600
rect 6886 27560 16574 27588
rect 18559 27560 18604 27588
rect 2222 27452 2228 27464
rect 2135 27424 2228 27452
rect 2222 27412 2228 27424
rect 2280 27452 2286 27464
rect 6886 27452 6914 27560
rect 9766 27520 9772 27532
rect 9727 27492 9772 27520
rect 9766 27480 9772 27492
rect 9824 27480 9830 27532
rect 9950 27480 9956 27532
rect 10008 27520 10014 27532
rect 10229 27523 10287 27529
rect 10229 27520 10241 27523
rect 10008 27492 10241 27520
rect 10008 27480 10014 27492
rect 10229 27489 10241 27492
rect 10275 27489 10287 27523
rect 16546 27520 16574 27560
rect 18598 27548 18604 27560
rect 18656 27548 18662 27600
rect 18782 27548 18788 27600
rect 18840 27588 18846 27600
rect 18840 27560 19564 27588
rect 18840 27548 18846 27560
rect 19426 27520 19432 27532
rect 16546 27492 19432 27520
rect 10229 27483 10287 27489
rect 19426 27480 19432 27492
rect 19484 27480 19490 27532
rect 19536 27529 19564 27560
rect 20070 27548 20076 27600
rect 20128 27588 20134 27600
rect 20622 27588 20628 27600
rect 20128 27560 20628 27588
rect 20128 27548 20134 27560
rect 20622 27548 20628 27560
rect 20680 27588 20686 27600
rect 28074 27588 28080 27600
rect 20680 27560 28080 27588
rect 20680 27548 20686 27560
rect 28074 27548 28080 27560
rect 28132 27548 28138 27600
rect 19521 27523 19579 27529
rect 19521 27489 19533 27523
rect 19567 27489 19579 27523
rect 19521 27483 19579 27489
rect 20993 27523 21051 27529
rect 20993 27489 21005 27523
rect 21039 27520 21051 27523
rect 21818 27520 21824 27532
rect 21039 27492 21824 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 21818 27480 21824 27492
rect 21876 27480 21882 27532
rect 22002 27520 22008 27532
rect 21963 27492 22008 27520
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 23290 27520 23296 27532
rect 23251 27492 23296 27520
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 9122 27452 9128 27464
rect 2280 27424 6914 27452
rect 9035 27424 9128 27452
rect 2280 27412 2286 27424
rect 9122 27412 9128 27424
rect 9180 27452 9186 27464
rect 9180 27424 9812 27452
rect 9180 27412 9186 27424
rect 9784 27316 9812 27424
rect 17402 27412 17408 27464
rect 17460 27452 17466 27464
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17460 27424 17601 27452
rect 17460 27412 17466 27424
rect 17589 27421 17601 27424
rect 17635 27452 17647 27455
rect 17862 27452 17868 27464
rect 17635 27424 17868 27452
rect 17635 27421 17647 27424
rect 17589 27415 17647 27421
rect 17862 27412 17868 27424
rect 17920 27412 17926 27464
rect 18322 27452 18328 27464
rect 18235 27424 18328 27452
rect 18322 27412 18328 27424
rect 18380 27452 18386 27464
rect 18782 27452 18788 27464
rect 18380 27424 18788 27452
rect 18380 27412 18386 27424
rect 18782 27412 18788 27424
rect 18840 27412 18846 27464
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27421 20867 27455
rect 22646 27452 22652 27464
rect 20809 27415 20867 27421
rect 21744 27424 22652 27452
rect 9950 27384 9956 27396
rect 9911 27356 9956 27384
rect 9950 27344 9956 27356
rect 10008 27344 10014 27396
rect 17880 27384 17908 27412
rect 19260 27384 19288 27415
rect 17880 27356 19288 27384
rect 20824 27384 20852 27415
rect 20824 27356 21496 27384
rect 10226 27316 10232 27328
rect 9784 27288 10232 27316
rect 10226 27276 10232 27288
rect 10284 27276 10290 27328
rect 17681 27319 17739 27325
rect 17681 27285 17693 27319
rect 17727 27316 17739 27319
rect 19334 27316 19340 27328
rect 17727 27288 19340 27316
rect 17727 27285 17739 27288
rect 17681 27279 17739 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 20346 27276 20352 27328
rect 20404 27316 20410 27328
rect 21468 27325 21496 27356
rect 21744 27328 21772 27424
rect 22646 27412 22652 27424
rect 22704 27412 22710 27464
rect 23014 27452 23020 27464
rect 22975 27424 23020 27452
rect 23014 27412 23020 27424
rect 23072 27412 23078 27464
rect 31754 27412 31760 27464
rect 31812 27452 31818 27464
rect 32677 27455 32735 27461
rect 32677 27452 32689 27455
rect 31812 27424 32689 27452
rect 31812 27412 31818 27424
rect 32677 27421 32689 27424
rect 32723 27421 32735 27455
rect 32677 27415 32735 27421
rect 21821 27387 21879 27393
rect 21821 27353 21833 27387
rect 21867 27384 21879 27387
rect 22462 27384 22468 27396
rect 21867 27356 22468 27384
rect 21867 27353 21879 27356
rect 21821 27347 21879 27353
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 20625 27319 20683 27325
rect 20625 27316 20637 27319
rect 20404 27288 20637 27316
rect 20404 27276 20410 27288
rect 20625 27285 20637 27288
rect 20671 27285 20683 27319
rect 20625 27279 20683 27285
rect 21453 27319 21511 27325
rect 21453 27285 21465 27319
rect 21499 27285 21511 27319
rect 21453 27279 21511 27285
rect 21726 27276 21732 27328
rect 21784 27316 21790 27328
rect 21913 27319 21971 27325
rect 21913 27316 21925 27319
rect 21784 27288 21925 27316
rect 21784 27276 21790 27288
rect 21913 27285 21925 27288
rect 21959 27285 21971 27319
rect 21913 27279 21971 27285
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 22649 27319 22707 27325
rect 22649 27316 22661 27319
rect 22336 27288 22661 27316
rect 22336 27276 22342 27288
rect 22649 27285 22661 27288
rect 22695 27285 22707 27319
rect 22649 27279 22707 27285
rect 22922 27276 22928 27328
rect 22980 27316 22986 27328
rect 23109 27319 23167 27325
rect 23109 27316 23121 27319
rect 22980 27288 23121 27316
rect 22980 27276 22986 27288
rect 23109 27285 23121 27288
rect 23155 27285 23167 27319
rect 23109 27279 23167 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 9950 27112 9956 27124
rect 9911 27084 9956 27112
rect 9950 27072 9956 27084
rect 10008 27072 10014 27124
rect 10226 27072 10232 27124
rect 10284 27112 10290 27124
rect 19426 27112 19432 27124
rect 10284 27084 19432 27112
rect 10284 27072 10290 27084
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 21821 27115 21879 27121
rect 21821 27112 21833 27115
rect 21600 27084 21833 27112
rect 21600 27072 21606 27084
rect 21821 27081 21833 27084
rect 21867 27081 21879 27115
rect 21821 27075 21879 27081
rect 22189 27115 22247 27121
rect 22189 27081 22201 27115
rect 22235 27112 22247 27115
rect 23014 27112 23020 27124
rect 22235 27084 23020 27112
rect 22235 27081 22247 27084
rect 22189 27075 22247 27081
rect 23014 27072 23020 27084
rect 23072 27072 23078 27124
rect 18601 27047 18659 27053
rect 18601 27044 18613 27047
rect 9876 27016 18613 27044
rect 9876 26985 9904 27016
rect 18601 27013 18613 27016
rect 18647 27044 18659 27047
rect 18690 27044 18696 27056
rect 18647 27016 18696 27044
rect 18647 27013 18659 27016
rect 18601 27007 18659 27013
rect 18690 27004 18696 27016
rect 18748 27004 18754 27056
rect 20070 27044 20076 27056
rect 20031 27016 20076 27044
rect 20070 27004 20076 27016
rect 20128 27004 20134 27056
rect 20806 27004 20812 27056
rect 20864 27044 20870 27056
rect 20993 27047 21051 27053
rect 20993 27044 21005 27047
rect 20864 27016 21005 27044
rect 20864 27004 20870 27016
rect 20993 27013 21005 27016
rect 21039 27013 21051 27047
rect 20993 27007 21051 27013
rect 22066 27016 31754 27044
rect 9861 26979 9919 26985
rect 9861 26945 9873 26979
rect 9907 26945 9919 26979
rect 9861 26939 9919 26945
rect 15194 26936 15200 26988
rect 15252 26976 15258 26988
rect 17405 26979 17463 26985
rect 15252 26974 16528 26976
rect 16592 26974 17172 26976
rect 15252 26948 17172 26974
rect 15252 26936 15258 26948
rect 16500 26946 16620 26948
rect 17144 26840 17172 26948
rect 17405 26945 17417 26979
rect 17451 26976 17463 26979
rect 17865 26979 17923 26985
rect 17865 26976 17877 26979
rect 17451 26948 17877 26976
rect 17451 26945 17463 26948
rect 17405 26939 17463 26945
rect 17865 26945 17877 26948
rect 17911 26976 17923 26979
rect 18322 26976 18328 26988
rect 17911 26948 18328 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 19334 26976 19340 26988
rect 19295 26948 19340 26976
rect 19334 26936 19340 26948
rect 19392 26976 19398 26988
rect 20530 26976 20536 26988
rect 19392 26948 20536 26976
rect 19392 26936 19398 26948
rect 20530 26936 20536 26948
rect 20588 26976 20594 26988
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 20588 26948 20729 26976
rect 20588 26936 20594 26948
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 21008 26976 21036 27007
rect 22066 26976 22094 27016
rect 21008 26948 22094 26976
rect 22281 26979 22339 26985
rect 20717 26939 20775 26945
rect 22281 26945 22293 26979
rect 22327 26976 22339 26979
rect 22922 26976 22928 26988
rect 22327 26948 22928 26976
rect 22327 26945 22339 26948
rect 22281 26939 22339 26945
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 22373 26911 22431 26917
rect 17276 26880 17321 26908
rect 17276 26868 17282 26880
rect 22373 26877 22385 26911
rect 22419 26877 22431 26911
rect 22373 26871 22431 26877
rect 22002 26840 22008 26852
rect 17144 26812 22008 26840
rect 22002 26800 22008 26812
rect 22060 26840 22066 26852
rect 22388 26840 22416 26871
rect 22060 26812 22416 26840
rect 22060 26800 22066 26812
rect 10778 26732 10784 26784
rect 10836 26772 10842 26784
rect 20070 26772 20076 26784
rect 10836 26744 20076 26772
rect 10836 26732 10842 26744
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 22370 26732 22376 26784
rect 22428 26772 22434 26784
rect 22480 26772 22508 26948
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 23198 26976 23204 26988
rect 23159 26948 23204 26976
rect 23198 26936 23204 26948
rect 23256 26936 23262 26988
rect 23382 26908 23388 26920
rect 23343 26880 23388 26908
rect 23382 26868 23388 26880
rect 23440 26868 23446 26920
rect 31726 26908 31754 27016
rect 38010 26976 38016 26988
rect 37971 26948 38016 26976
rect 38010 26936 38016 26948
rect 38068 26936 38074 26988
rect 37274 26908 37280 26920
rect 31726 26880 37280 26908
rect 37274 26868 37280 26880
rect 37332 26868 37338 26920
rect 22428 26744 22508 26772
rect 22428 26732 22434 26744
rect 22554 26732 22560 26784
rect 22612 26772 22618 26784
rect 23017 26775 23075 26781
rect 23017 26772 23029 26775
rect 22612 26744 23029 26772
rect 22612 26732 22618 26744
rect 23017 26741 23029 26744
rect 23063 26772 23075 26775
rect 23198 26772 23204 26784
rect 23063 26744 23204 26772
rect 23063 26741 23075 26744
rect 23017 26735 23075 26741
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 23842 26732 23848 26784
rect 23900 26772 23906 26784
rect 37921 26775 37979 26781
rect 37921 26772 37933 26775
rect 23900 26744 37933 26772
rect 23900 26732 23906 26744
rect 37921 26741 37933 26744
rect 37967 26741 37979 26775
rect 37921 26735 37979 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 18230 26528 18236 26580
rect 18288 26568 18294 26580
rect 28074 26568 28080 26580
rect 18288 26540 28080 26568
rect 18288 26528 18294 26540
rect 28074 26528 28080 26540
rect 28132 26528 28138 26580
rect 6886 26472 22094 26500
rect 2038 26392 2044 26444
rect 2096 26432 2102 26444
rect 6886 26432 6914 26472
rect 18230 26432 18236 26444
rect 2096 26404 6914 26432
rect 18191 26404 18236 26432
rect 2096 26392 2102 26404
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 19426 26392 19432 26444
rect 19484 26432 19490 26444
rect 19705 26435 19763 26441
rect 19705 26432 19717 26435
rect 19484 26404 19717 26432
rect 19484 26392 19490 26404
rect 19705 26401 19717 26404
rect 19751 26432 19763 26435
rect 19978 26432 19984 26444
rect 19751 26404 19984 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 19978 26392 19984 26404
rect 20036 26392 20042 26444
rect 22066 26432 22094 26472
rect 22066 26404 23428 26432
rect 1578 26324 1584 26376
rect 1636 26364 1642 26376
rect 1673 26367 1731 26373
rect 1673 26364 1685 26367
rect 1636 26336 1685 26364
rect 1636 26324 1642 26336
rect 1673 26333 1685 26336
rect 1719 26333 1731 26367
rect 17494 26364 17500 26376
rect 17455 26336 17500 26364
rect 1673 26327 1731 26333
rect 17494 26324 17500 26336
rect 17552 26324 17558 26376
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 18601 26367 18659 26373
rect 18601 26364 18613 26367
rect 18380 26336 18613 26364
rect 18380 26324 18386 26336
rect 18601 26333 18613 26336
rect 18647 26333 18659 26367
rect 20530 26364 20536 26376
rect 20491 26336 20536 26364
rect 18601 26327 18659 26333
rect 20530 26324 20536 26336
rect 20588 26324 20594 26376
rect 21174 26324 21180 26376
rect 21232 26364 21238 26376
rect 22112 26373 22140 26404
rect 23400 26376 23428 26404
rect 21269 26367 21327 26373
rect 21269 26364 21281 26367
rect 21232 26336 21281 26364
rect 21232 26324 21238 26336
rect 21269 26333 21281 26336
rect 21315 26333 21327 26367
rect 21269 26327 21327 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22278 26364 22284 26376
rect 22239 26336 22284 26364
rect 22097 26327 22155 26333
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 22554 26364 22560 26376
rect 22515 26336 22560 26364
rect 22554 26324 22560 26336
rect 22612 26324 22618 26376
rect 22738 26364 22744 26376
rect 22699 26336 22744 26364
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23382 26364 23388 26376
rect 23343 26336 23388 26364
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 34698 26364 34704 26376
rect 34659 26336 34704 26364
rect 34698 26324 34704 26336
rect 34756 26324 34762 26376
rect 36262 26364 36268 26376
rect 36223 26336 36268 26364
rect 36262 26324 36268 26336
rect 36320 26324 36326 26376
rect 21082 26296 21088 26308
rect 21043 26268 21088 26296
rect 21082 26256 21088 26268
rect 21140 26256 21146 26308
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 21453 26299 21511 26305
rect 21453 26296 21465 26299
rect 21416 26268 21465 26296
rect 21416 26256 21422 26268
rect 21453 26265 21465 26268
rect 21499 26265 21511 26299
rect 22296 26296 22324 26324
rect 23201 26299 23259 26305
rect 23201 26296 23213 26299
rect 22296 26268 23213 26296
rect 21453 26259 21511 26265
rect 23201 26265 23213 26268
rect 23247 26265 23259 26299
rect 23201 26259 23259 26265
rect 23290 26256 23296 26308
rect 23348 26296 23354 26308
rect 23569 26299 23627 26305
rect 23569 26296 23581 26299
rect 23348 26268 23581 26296
rect 23348 26256 23354 26268
rect 23569 26265 23581 26268
rect 23615 26265 23627 26299
rect 23569 26259 23627 26265
rect 36449 26299 36507 26305
rect 36449 26265 36461 26299
rect 36495 26296 36507 26299
rect 37366 26296 37372 26308
rect 36495 26268 37372 26296
rect 36495 26265 36507 26268
rect 36449 26259 36507 26265
rect 37366 26256 37372 26268
rect 37424 26256 37430 26308
rect 38105 26299 38163 26305
rect 38105 26265 38117 26299
rect 38151 26296 38163 26299
rect 38194 26296 38200 26308
rect 38151 26268 38200 26296
rect 38151 26265 38163 26268
rect 38105 26259 38163 26265
rect 38194 26256 38200 26268
rect 38252 26256 38258 26308
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 22186 25984 22192 26036
rect 22244 26024 22250 26036
rect 22833 26027 22891 26033
rect 22833 26024 22845 26027
rect 22244 25996 22845 26024
rect 22244 25984 22250 25996
rect 22833 25993 22845 25996
rect 22879 26024 22891 26027
rect 23014 26024 23020 26036
rect 22879 25996 23020 26024
rect 22879 25993 22891 25996
rect 22833 25987 22891 25993
rect 23014 25984 23020 25996
rect 23072 25984 23078 26036
rect 23201 26027 23259 26033
rect 23201 25993 23213 26027
rect 23247 26024 23259 26027
rect 23382 26024 23388 26036
rect 23247 25996 23388 26024
rect 23247 25993 23259 25996
rect 23201 25987 23259 25993
rect 23382 25984 23388 25996
rect 23440 26024 23446 26036
rect 37366 26024 37372 26036
rect 23440 25996 23704 26024
rect 37327 25996 37372 26024
rect 23440 25984 23446 25996
rect 3418 25956 3424 25968
rect 3379 25928 3424 25956
rect 3418 25916 3424 25928
rect 3476 25916 3482 25968
rect 18414 25956 18420 25968
rect 17144 25928 18420 25956
rect 17144 25900 17172 25928
rect 18414 25916 18420 25928
rect 18472 25916 18478 25968
rect 23676 25965 23704 25996
rect 37366 25984 37372 25996
rect 37424 25984 37430 26036
rect 23661 25959 23719 25965
rect 23661 25925 23673 25959
rect 23707 25925 23719 25959
rect 23842 25956 23848 25968
rect 23803 25928 23848 25956
rect 23661 25919 23719 25925
rect 23842 25916 23848 25928
rect 23900 25916 23906 25968
rect 33505 25959 33563 25965
rect 33505 25925 33517 25959
rect 33551 25956 33563 25959
rect 34241 25959 34299 25965
rect 34241 25956 34253 25959
rect 33551 25928 34253 25956
rect 33551 25925 33563 25928
rect 33505 25919 33563 25925
rect 34241 25925 34253 25928
rect 34287 25925 34299 25959
rect 34241 25919 34299 25925
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 17126 25888 17132 25900
rect 17087 25860 17132 25888
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 17494 25848 17500 25900
rect 17552 25888 17558 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17552 25860 17601 25888
rect 17552 25848 17558 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 20530 25888 20536 25900
rect 20491 25860 20536 25888
rect 17589 25851 17647 25857
rect 20530 25848 20536 25860
rect 20588 25848 20594 25900
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21232 25860 21833 25888
rect 21232 25848 21238 25860
rect 21821 25857 21833 25860
rect 21867 25888 21879 25891
rect 21910 25888 21916 25900
rect 21867 25860 21916 25888
rect 21867 25857 21879 25860
rect 21821 25851 21879 25857
rect 21910 25848 21916 25860
rect 21968 25848 21974 25900
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25888 22063 25891
rect 22094 25888 22100 25900
rect 22051 25860 22100 25888
rect 22051 25857 22063 25860
rect 22005 25851 22063 25857
rect 22094 25848 22100 25860
rect 22152 25848 22158 25900
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 22741 25891 22799 25897
rect 22741 25888 22753 25891
rect 22428 25860 22753 25888
rect 22428 25848 22434 25860
rect 22741 25857 22753 25860
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 33318 25848 33324 25900
rect 33376 25888 33382 25900
rect 33413 25891 33471 25897
rect 33413 25888 33425 25891
rect 33376 25860 33425 25888
rect 33376 25848 33382 25860
rect 33413 25857 33425 25860
rect 33459 25857 33471 25891
rect 33413 25851 33471 25857
rect 36262 25848 36268 25900
rect 36320 25888 36326 25900
rect 36541 25891 36599 25897
rect 36541 25888 36553 25891
rect 36320 25860 36553 25888
rect 36320 25848 36326 25860
rect 36541 25857 36553 25860
rect 36587 25857 36599 25891
rect 37274 25888 37280 25900
rect 37235 25860 37280 25888
rect 36541 25851 36599 25857
rect 37274 25848 37280 25860
rect 37332 25848 37338 25900
rect 37918 25888 37924 25900
rect 37879 25860 37924 25888
rect 37918 25848 37924 25860
rect 37976 25848 37982 25900
rect 1765 25823 1823 25829
rect 1765 25789 1777 25823
rect 1811 25820 1823 25823
rect 2038 25820 2044 25832
rect 1811 25792 2044 25820
rect 1811 25789 1823 25792
rect 1765 25783 1823 25789
rect 2038 25780 2044 25792
rect 2096 25780 2102 25832
rect 3510 25780 3516 25832
rect 3568 25820 3574 25832
rect 17037 25823 17095 25829
rect 3568 25792 6914 25820
rect 3568 25780 3574 25792
rect 6886 25752 6914 25792
rect 17037 25789 17049 25823
rect 17083 25820 17095 25823
rect 17773 25823 17831 25829
rect 17773 25820 17785 25823
rect 17083 25792 17785 25820
rect 17083 25789 17095 25792
rect 17037 25783 17095 25789
rect 17773 25789 17785 25792
rect 17819 25789 17831 25823
rect 17773 25783 17831 25789
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 20257 25823 20315 25829
rect 20257 25789 20269 25823
rect 20303 25820 20315 25823
rect 20438 25820 20444 25832
rect 20303 25792 20444 25820
rect 20303 25789 20315 25792
rect 20257 25783 20315 25789
rect 18064 25752 18092 25783
rect 20438 25780 20444 25792
rect 20496 25780 20502 25832
rect 22646 25820 22652 25832
rect 22607 25792 22652 25820
rect 22646 25780 22652 25792
rect 22704 25780 22710 25832
rect 34057 25823 34115 25829
rect 34057 25789 34069 25823
rect 34103 25820 34115 25823
rect 34698 25820 34704 25832
rect 34103 25792 34704 25820
rect 34103 25789 34115 25792
rect 34057 25783 34115 25789
rect 34698 25780 34704 25792
rect 34756 25780 34762 25832
rect 35802 25820 35808 25832
rect 35763 25792 35808 25820
rect 35802 25780 35808 25792
rect 35860 25780 35866 25832
rect 6886 25724 18092 25752
rect 20456 25752 20484 25780
rect 37458 25752 37464 25764
rect 20456 25724 37464 25752
rect 37458 25712 37464 25724
rect 37516 25712 37522 25764
rect 21913 25687 21971 25693
rect 21913 25653 21925 25687
rect 21959 25684 21971 25687
rect 23474 25684 23480 25696
rect 21959 25656 23480 25684
rect 21959 25653 21971 25656
rect 21913 25647 21971 25653
rect 23474 25644 23480 25656
rect 23532 25644 23538 25696
rect 24026 25684 24032 25696
rect 23987 25656 24032 25684
rect 24026 25644 24032 25656
rect 24084 25644 24090 25696
rect 37918 25644 37924 25696
rect 37976 25684 37982 25696
rect 38013 25687 38071 25693
rect 38013 25684 38025 25687
rect 37976 25656 38025 25684
rect 37976 25644 37982 25656
rect 38013 25653 38025 25656
rect 38059 25653 38071 25687
rect 38013 25647 38071 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2038 25480 2044 25492
rect 1999 25452 2044 25480
rect 2038 25440 2044 25452
rect 2096 25440 2102 25492
rect 20717 25483 20775 25489
rect 20717 25449 20729 25483
rect 20763 25480 20775 25483
rect 21082 25480 21088 25492
rect 20763 25452 21088 25480
rect 20763 25449 20775 25452
rect 20717 25443 20775 25449
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 21542 25440 21548 25492
rect 21600 25480 21606 25492
rect 22462 25480 22468 25492
rect 21600 25452 22468 25480
rect 21600 25440 21606 25452
rect 22462 25440 22468 25452
rect 22520 25440 22526 25492
rect 22646 25480 22652 25492
rect 22559 25452 22652 25480
rect 22370 25412 22376 25424
rect 19904 25384 22376 25412
rect 2133 25279 2191 25285
rect 2133 25245 2145 25279
rect 2179 25276 2191 25279
rect 2314 25276 2320 25288
rect 2179 25248 2320 25276
rect 2179 25245 2191 25248
rect 2133 25239 2191 25245
rect 2314 25236 2320 25248
rect 2372 25276 2378 25288
rect 18598 25276 18604 25288
rect 2372 25248 6914 25276
rect 18559 25248 18604 25276
rect 2372 25236 2378 25248
rect 6886 25208 6914 25248
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 19904 25276 19932 25384
rect 22370 25372 22376 25384
rect 22428 25372 22434 25424
rect 20070 25344 20076 25356
rect 20031 25316 20076 25344
rect 20070 25304 20076 25316
rect 20128 25344 20134 25356
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 20128 25316 21281 25344
rect 20128 25304 20134 25316
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 21269 25307 21327 25313
rect 21453 25347 21511 25353
rect 21453 25313 21465 25347
rect 21499 25344 21511 25347
rect 21726 25344 21732 25356
rect 21499 25316 21732 25344
rect 21499 25313 21511 25316
rect 21453 25307 21511 25313
rect 21726 25304 21732 25316
rect 21784 25344 21790 25356
rect 21784 25316 22416 25344
rect 21784 25304 21790 25316
rect 20257 25279 20315 25285
rect 20257 25276 20269 25279
rect 19904 25248 20269 25276
rect 20257 25245 20269 25248
rect 20303 25245 20315 25279
rect 20257 25239 20315 25245
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25276 20407 25279
rect 22186 25276 22192 25288
rect 20395 25248 22192 25276
rect 20395 25245 20407 25248
rect 20349 25239 20407 25245
rect 22186 25236 22192 25248
rect 22244 25236 22250 25288
rect 17954 25208 17960 25220
rect 6886 25180 17960 25208
rect 17954 25168 17960 25180
rect 18012 25208 18018 25220
rect 18049 25211 18107 25217
rect 18049 25208 18061 25211
rect 18012 25180 18061 25208
rect 18012 25168 18018 25180
rect 18049 25177 18061 25180
rect 18095 25177 18107 25211
rect 21542 25208 21548 25220
rect 21503 25180 21548 25208
rect 18049 25171 18107 25177
rect 21542 25168 21548 25180
rect 21600 25168 21606 25220
rect 22388 25208 22416 25316
rect 22462 25304 22468 25356
rect 22520 25304 22526 25356
rect 22572 25353 22600 25452
rect 22646 25440 22652 25452
rect 22704 25480 22710 25492
rect 22704 25452 28994 25480
rect 22704 25440 22710 25452
rect 25225 25415 25283 25421
rect 25225 25381 25237 25415
rect 25271 25412 25283 25415
rect 28966 25412 28994 25452
rect 37826 25412 37832 25424
rect 25271 25384 25728 25412
rect 28966 25384 37832 25412
rect 25271 25381 25283 25384
rect 25225 25375 25283 25381
rect 25700 25353 25728 25384
rect 37826 25372 37832 25384
rect 37884 25372 37890 25424
rect 22557 25347 22615 25353
rect 22557 25313 22569 25347
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 25685 25347 25743 25353
rect 25685 25313 25697 25347
rect 25731 25313 25743 25347
rect 25685 25307 25743 25313
rect 27525 25347 27583 25353
rect 27525 25313 27537 25347
rect 27571 25344 27583 25347
rect 28258 25344 28264 25356
rect 27571 25316 28264 25344
rect 27571 25313 27583 25316
rect 27525 25307 27583 25313
rect 28258 25304 28264 25316
rect 28316 25304 28322 25356
rect 37918 25344 37924 25356
rect 37879 25316 37924 25344
rect 37918 25304 37924 25316
rect 37976 25304 37982 25356
rect 22480 25276 22508 25304
rect 22741 25279 22799 25285
rect 22741 25276 22753 25279
rect 22480 25248 22753 25276
rect 22741 25245 22753 25248
rect 22787 25245 22799 25279
rect 23569 25279 23627 25285
rect 23569 25276 23581 25279
rect 22741 25239 22799 25245
rect 23124 25248 23581 25276
rect 22388 25180 22600 25208
rect 22572 25152 22600 25180
rect 21913 25143 21971 25149
rect 21913 25109 21925 25143
rect 21959 25140 21971 25143
rect 22094 25140 22100 25152
rect 21959 25112 22100 25140
rect 21959 25109 21971 25112
rect 21913 25103 21971 25109
rect 22094 25100 22100 25112
rect 22152 25140 22158 25152
rect 22462 25140 22468 25152
rect 22152 25112 22468 25140
rect 22152 25100 22158 25112
rect 22462 25100 22468 25112
rect 22520 25100 22526 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22649 25143 22707 25149
rect 22649 25140 22661 25143
rect 22612 25112 22661 25140
rect 22612 25100 22618 25112
rect 22649 25109 22661 25112
rect 22695 25109 22707 25143
rect 22649 25103 22707 25109
rect 23014 25100 23020 25152
rect 23072 25140 23078 25152
rect 23124 25149 23152 25248
rect 23569 25245 23581 25248
rect 23615 25245 23627 25279
rect 23569 25239 23627 25245
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25276 23811 25279
rect 23842 25276 23848 25288
rect 23799 25248 23848 25276
rect 23799 25245 23811 25248
rect 23753 25239 23811 25245
rect 23842 25236 23848 25248
rect 23900 25236 23906 25288
rect 24302 25236 24308 25288
rect 24360 25276 24366 25288
rect 25041 25279 25099 25285
rect 25041 25276 25053 25279
rect 24360 25248 25053 25276
rect 24360 25236 24366 25248
rect 25041 25245 25053 25248
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 38102 25236 38108 25288
rect 38160 25276 38166 25288
rect 38160 25248 38205 25276
rect 38160 25236 38166 25248
rect 25866 25208 25872 25220
rect 25827 25180 25872 25208
rect 25866 25168 25872 25180
rect 25924 25168 25930 25220
rect 36170 25168 36176 25220
rect 36228 25208 36234 25220
rect 36265 25211 36323 25217
rect 36265 25208 36277 25211
rect 36228 25180 36277 25208
rect 36228 25168 36234 25180
rect 36265 25177 36277 25180
rect 36311 25177 36323 25211
rect 36265 25171 36323 25177
rect 23109 25143 23167 25149
rect 23109 25140 23121 25143
rect 23072 25112 23121 25140
rect 23072 25100 23078 25112
rect 23109 25109 23121 25112
rect 23155 25109 23167 25143
rect 23109 25103 23167 25109
rect 23566 25100 23572 25152
rect 23624 25140 23630 25152
rect 23661 25143 23719 25149
rect 23661 25140 23673 25143
rect 23624 25112 23673 25140
rect 23624 25100 23630 25112
rect 23661 25109 23673 25112
rect 23707 25109 23719 25143
rect 23661 25103 23719 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 24302 24936 24308 24948
rect 22204 24908 23520 24936
rect 24263 24908 24308 24936
rect 22204 24877 22232 24908
rect 22189 24871 22247 24877
rect 22189 24837 22201 24871
rect 22235 24837 22247 24871
rect 23014 24868 23020 24880
rect 22189 24831 22247 24837
rect 22301 24840 23020 24868
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24800 18475 24803
rect 18598 24800 18604 24812
rect 18463 24772 18604 24800
rect 18463 24769 18475 24772
rect 18417 24763 18475 24769
rect 18598 24760 18604 24772
rect 18656 24800 18662 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 18656 24772 19717 24800
rect 18656 24760 18662 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 20530 24800 20536 24812
rect 20491 24772 20536 24800
rect 19705 24763 19763 24769
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 21082 24760 21088 24812
rect 21140 24800 21146 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21140 24772 21833 24800
rect 21140 24760 21146 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 21910 24760 21916 24812
rect 21968 24800 21974 24812
rect 22094 24809 22100 24812
rect 22051 24803 22100 24809
rect 21968 24772 22013 24800
rect 21968 24760 21974 24772
rect 22051 24769 22063 24803
rect 22097 24769 22100 24803
rect 22051 24763 22100 24769
rect 22094 24760 22100 24763
rect 22152 24760 22158 24812
rect 22301 24809 22329 24840
rect 23014 24828 23020 24840
rect 23072 24828 23078 24880
rect 22301 24803 22363 24809
rect 22301 24772 22317 24803
rect 22305 24769 22317 24772
rect 22351 24769 22363 24803
rect 22305 24763 22363 24769
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 23109 24803 23167 24809
rect 23109 24800 23121 24803
rect 22520 24772 23121 24800
rect 22520 24760 22526 24772
rect 23109 24769 23121 24772
rect 23155 24769 23167 24803
rect 23109 24763 23167 24769
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23382 24800 23388 24812
rect 23343 24772 23388 24800
rect 23201 24763 23259 24769
rect 19058 24732 19064 24744
rect 19019 24704 19064 24732
rect 19058 24692 19064 24704
rect 19116 24692 19122 24744
rect 4798 24624 4804 24676
rect 4856 24664 4862 24676
rect 20548 24664 20576 24760
rect 21929 24732 21957 24760
rect 23216 24732 23244 24763
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 23492 24809 23520 24908
rect 24302 24896 24308 24908
rect 24360 24896 24366 24948
rect 25866 24936 25872 24948
rect 25827 24908 25872 24936
rect 25866 24896 25872 24908
rect 25924 24896 25930 24948
rect 23566 24828 23572 24880
rect 23624 24868 23630 24880
rect 23624 24840 24808 24868
rect 23624 24828 23630 24840
rect 23477 24803 23535 24809
rect 23477 24769 23489 24803
rect 23523 24800 23535 24803
rect 23842 24800 23848 24812
rect 23523 24772 23848 24800
rect 23523 24769 23535 24772
rect 23477 24763 23535 24769
rect 23842 24760 23848 24772
rect 23900 24760 23906 24812
rect 24780 24809 24808 24840
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24769 23995 24803
rect 23937 24763 23995 24769
rect 24765 24803 24823 24809
rect 24765 24769 24777 24803
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 24949 24763 25007 24769
rect 23952 24732 23980 24763
rect 21929 24704 23244 24732
rect 23584 24704 23980 24732
rect 24029 24735 24087 24741
rect 4856 24636 20576 24664
rect 4856 24624 4862 24636
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 22925 24667 22983 24673
rect 22925 24664 22937 24667
rect 21324 24636 22937 24664
rect 21324 24624 21330 24636
rect 22925 24633 22937 24636
rect 22971 24664 22983 24667
rect 23382 24664 23388 24676
rect 22971 24636 23388 24664
rect 22971 24633 22983 24636
rect 22925 24627 22983 24633
rect 23382 24624 23388 24636
rect 23440 24624 23446 24676
rect 19058 24556 19064 24608
rect 19116 24596 19122 24608
rect 21450 24596 21456 24608
rect 19116 24568 21456 24596
rect 19116 24556 19122 24568
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 22465 24599 22523 24605
rect 22465 24596 22477 24599
rect 21968 24568 22477 24596
rect 21968 24556 21974 24568
rect 22465 24565 22477 24568
rect 22511 24565 22523 24599
rect 22465 24559 22523 24565
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 23584 24596 23612 24704
rect 24029 24701 24041 24735
rect 24075 24732 24087 24735
rect 24857 24735 24915 24741
rect 24857 24732 24869 24735
rect 24075 24704 24869 24732
rect 24075 24701 24087 24704
rect 24029 24695 24087 24701
rect 24857 24701 24869 24704
rect 24903 24701 24915 24735
rect 24857 24695 24915 24701
rect 23750 24624 23756 24676
rect 23808 24664 23814 24676
rect 24964 24664 24992 24763
rect 25590 24760 25596 24812
rect 25648 24800 25654 24812
rect 25777 24803 25835 24809
rect 25777 24800 25789 24803
rect 25648 24772 25789 24800
rect 25648 24760 25654 24772
rect 25777 24769 25789 24772
rect 25823 24769 25835 24803
rect 25777 24763 25835 24769
rect 37829 24803 37887 24809
rect 37829 24769 37841 24803
rect 37875 24800 37887 24803
rect 38102 24800 38108 24812
rect 37875 24772 38108 24800
rect 37875 24769 37887 24772
rect 37829 24763 37887 24769
rect 38102 24760 38108 24772
rect 38160 24760 38166 24812
rect 23808 24636 24992 24664
rect 23808 24624 23814 24636
rect 23256 24568 23612 24596
rect 23256 24556 23262 24568
rect 23658 24556 23664 24608
rect 23716 24596 23722 24608
rect 23937 24599 23995 24605
rect 23937 24596 23949 24599
rect 23716 24568 23949 24596
rect 23716 24556 23722 24568
rect 23937 24565 23949 24568
rect 23983 24565 23995 24599
rect 23937 24559 23995 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 21358 24392 21364 24404
rect 21008 24364 21364 24392
rect 17405 24327 17463 24333
rect 17405 24293 17417 24327
rect 17451 24324 17463 24327
rect 17451 24296 18092 24324
rect 17451 24293 17463 24296
rect 17405 24287 17463 24293
rect 18064 24256 18092 24296
rect 18598 24256 18604 24268
rect 18064 24228 18604 24256
rect 1854 24148 1860 24200
rect 1912 24188 1918 24200
rect 1949 24191 2007 24197
rect 1949 24188 1961 24191
rect 1912 24160 1961 24188
rect 1912 24148 1918 24160
rect 1949 24157 1961 24160
rect 1995 24157 2007 24191
rect 17218 24188 17224 24200
rect 17179 24160 17224 24188
rect 1949 24151 2007 24157
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 18064 24197 18092 24228
rect 18598 24216 18604 24228
rect 18656 24216 18662 24268
rect 21008 24256 21036 24364
rect 21358 24352 21364 24364
rect 21416 24392 21422 24404
rect 22554 24392 22560 24404
rect 21416 24364 22560 24392
rect 21416 24352 21422 24364
rect 22554 24352 22560 24364
rect 22612 24392 22618 24404
rect 22612 24364 23704 24392
rect 22612 24352 22618 24364
rect 21910 24324 21916 24336
rect 21192 24296 21916 24324
rect 21192 24265 21220 24296
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 22005 24327 22063 24333
rect 22005 24293 22017 24327
rect 22051 24324 22063 24327
rect 22830 24324 22836 24336
rect 22051 24296 22836 24324
rect 22051 24293 22063 24296
rect 22005 24287 22063 24293
rect 22830 24284 22836 24296
rect 22888 24284 22894 24336
rect 21085 24259 21143 24265
rect 21085 24256 21097 24259
rect 20180 24228 21097 24256
rect 20180 24197 20208 24228
rect 21085 24225 21097 24228
rect 21131 24225 21143 24259
rect 21085 24219 21143 24225
rect 21177 24259 21235 24265
rect 21177 24225 21189 24259
rect 21223 24225 21235 24259
rect 21928 24256 21956 24284
rect 21928 24228 23336 24256
rect 21177 24219 21235 24225
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24157 18107 24191
rect 18049 24151 18107 24157
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24157 20223 24191
rect 20346 24188 20352 24200
rect 20307 24160 20352 24188
rect 20165 24151 20223 24157
rect 18601 24123 18659 24129
rect 18601 24089 18613 24123
rect 18647 24120 18659 24123
rect 18782 24120 18788 24132
rect 18647 24092 18788 24120
rect 18647 24089 18659 24092
rect 18601 24083 18659 24089
rect 18782 24080 18788 24092
rect 18840 24080 18846 24132
rect 20088 24120 20116 24151
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 20441 24191 20499 24197
rect 20441 24157 20453 24191
rect 20487 24188 20499 24191
rect 20530 24188 20536 24200
rect 20487 24160 20536 24188
rect 20487 24157 20499 24160
rect 20441 24151 20499 24157
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20956 24160 21005 24188
rect 20956 24148 20962 24160
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 21266 24188 21272 24200
rect 21179 24160 21272 24188
rect 20993 24151 21051 24157
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 21284 24120 21312 24148
rect 20088 24092 21312 24120
rect 22020 24120 22048 24151
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 22189 24191 22247 24197
rect 22189 24188 22201 24191
rect 22152 24160 22201 24188
rect 22152 24148 22158 24160
rect 22189 24157 22201 24160
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 22572 24120 22600 24151
rect 22646 24148 22652 24200
rect 22704 24188 22710 24200
rect 22741 24191 22799 24197
rect 22741 24188 22753 24191
rect 22704 24160 22753 24188
rect 22704 24148 22710 24160
rect 22741 24157 22753 24160
rect 22787 24188 22799 24191
rect 23198 24188 23204 24200
rect 22787 24160 23204 24188
rect 22787 24157 22799 24160
rect 22741 24151 22799 24157
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 23308 24188 23336 24228
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 23569 24259 23627 24265
rect 23440 24228 23485 24256
rect 23440 24216 23446 24228
rect 23569 24225 23581 24259
rect 23615 24256 23627 24259
rect 23676 24256 23704 24364
rect 24394 24324 24400 24336
rect 24355 24296 24400 24324
rect 24394 24284 24400 24296
rect 24452 24284 24458 24336
rect 25498 24256 25504 24268
rect 23615 24228 23704 24256
rect 25459 24228 25504 24256
rect 23615 24225 23627 24228
rect 23569 24219 23627 24225
rect 25498 24216 25504 24228
rect 25556 24216 25562 24268
rect 27338 24256 27344 24268
rect 27299 24228 27344 24256
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 23477 24191 23535 24197
rect 23477 24188 23489 24191
rect 23308 24160 23489 24188
rect 23477 24157 23489 24160
rect 23523 24157 23535 24191
rect 23658 24188 23664 24200
rect 23619 24160 23664 24188
rect 23477 24151 23535 24157
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 24673 24191 24731 24197
rect 24673 24188 24685 24191
rect 23768 24160 24685 24188
rect 22020 24092 22094 24120
rect 22572 24092 23244 24120
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 21358 24052 21364 24064
rect 19935 24024 21364 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 21358 24012 21364 24024
rect 21416 24012 21422 24064
rect 21453 24055 21511 24061
rect 21453 24021 21465 24055
rect 21499 24052 21511 24055
rect 21818 24052 21824 24064
rect 21499 24024 21824 24052
rect 21499 24021 21511 24024
rect 21453 24015 21511 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22066 24052 22094 24092
rect 23106 24052 23112 24064
rect 22066 24024 23112 24052
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 23216 24061 23244 24092
rect 23290 24080 23296 24132
rect 23348 24120 23354 24132
rect 23676 24120 23704 24148
rect 23348 24092 23704 24120
rect 23348 24080 23354 24092
rect 23201 24055 23259 24061
rect 23201 24021 23213 24055
rect 23247 24052 23259 24055
rect 23768 24052 23796 24160
rect 24673 24157 24685 24160
rect 24719 24157 24731 24191
rect 24673 24151 24731 24157
rect 37829 24191 37887 24197
rect 37829 24157 37841 24191
rect 37875 24188 37887 24191
rect 38102 24188 38108 24200
rect 37875 24160 38108 24188
rect 37875 24157 37887 24160
rect 37829 24151 37887 24157
rect 38102 24148 38108 24160
rect 38160 24148 38166 24200
rect 23842 24080 23848 24132
rect 23900 24120 23906 24132
rect 24397 24123 24455 24129
rect 24397 24120 24409 24123
rect 23900 24092 24409 24120
rect 23900 24080 23906 24092
rect 24397 24089 24409 24092
rect 24443 24089 24455 24123
rect 25682 24120 25688 24132
rect 25643 24092 25688 24120
rect 24397 24083 24455 24089
rect 25682 24080 25688 24092
rect 25740 24080 25746 24132
rect 24578 24052 24584 24064
rect 23247 24024 23796 24052
rect 24539 24024 24584 24052
rect 23247 24021 23259 24024
rect 23201 24015 23259 24021
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 21082 23848 21088 23860
rect 21043 23820 21088 23848
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 25682 23848 25688 23860
rect 21416 23820 22324 23848
rect 25643 23820 25688 23848
rect 21416 23808 21422 23820
rect 3694 23780 3700 23792
rect 3655 23752 3700 23780
rect 3694 23740 3700 23752
rect 3752 23740 3758 23792
rect 18414 23780 18420 23792
rect 18375 23752 18420 23780
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 17218 23672 17224 23724
rect 17276 23712 17282 23724
rect 17862 23712 17868 23724
rect 17276 23684 17868 23712
rect 17276 23672 17282 23684
rect 17862 23672 17868 23684
rect 17920 23712 17926 23724
rect 17920 23684 18552 23712
rect 17920 23672 17926 23684
rect 2038 23644 2044 23656
rect 1999 23616 2044 23644
rect 2038 23604 2044 23616
rect 2096 23604 2102 23656
rect 18524 23644 18552 23684
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18656 23684 19073 23712
rect 18656 23672 18662 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19981 23715 20039 23721
rect 19981 23712 19993 23715
rect 19484 23684 19993 23712
rect 19484 23672 19490 23684
rect 19981 23681 19993 23684
rect 20027 23681 20039 23715
rect 20990 23712 20996 23724
rect 20951 23684 20996 23712
rect 19981 23675 20039 23681
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 22094 23712 22100 23724
rect 22055 23684 22100 23712
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 22186 23718 22244 23724
rect 22296 23721 22324 23820
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 22388 23752 22784 23780
rect 22186 23684 22198 23718
rect 22232 23684 22244 23718
rect 22186 23678 22244 23684
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 18524 23616 19717 23644
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 20530 23604 20536 23656
rect 20588 23644 20594 23656
rect 22204 23644 22232 23678
rect 22281 23675 22339 23681
rect 22388 23644 22416 23752
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23712 22523 23715
rect 22646 23712 22652 23724
rect 22511 23684 22652 23712
rect 22511 23681 22523 23684
rect 22465 23675 22523 23681
rect 22646 23672 22652 23684
rect 22704 23672 22710 23724
rect 22756 23712 22784 23752
rect 22830 23740 22836 23792
rect 22888 23780 22894 23792
rect 28166 23780 28172 23792
rect 22888 23752 28172 23780
rect 22888 23740 22894 23752
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 23106 23712 23112 23724
rect 22756 23684 23112 23712
rect 23106 23672 23112 23684
rect 23164 23672 23170 23724
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23712 23351 23715
rect 24394 23712 24400 23724
rect 23339 23684 24400 23712
rect 23339 23681 23351 23684
rect 23293 23675 23351 23681
rect 24394 23672 24400 23684
rect 24452 23672 24458 23724
rect 25590 23712 25596 23724
rect 25551 23684 25596 23712
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 37274 23712 37280 23724
rect 37235 23684 37280 23712
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 20588 23616 22416 23644
rect 20588 23604 20594 23616
rect 22738 23604 22744 23656
rect 22796 23644 22802 23656
rect 23201 23647 23259 23653
rect 23201 23644 23213 23647
rect 22796 23616 23213 23644
rect 22796 23604 22802 23616
rect 23201 23613 23213 23616
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 18598 23536 18604 23588
rect 18656 23576 18662 23588
rect 18782 23576 18788 23588
rect 18656 23548 18788 23576
rect 18656 23536 18662 23548
rect 18782 23536 18788 23548
rect 18840 23536 18846 23588
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 23290 23576 23296 23588
rect 20404 23548 23296 23576
rect 20404 23536 20410 23548
rect 23290 23536 23296 23548
rect 23348 23536 23354 23588
rect 21450 23468 21456 23520
rect 21508 23508 21514 23520
rect 21821 23511 21879 23517
rect 21821 23508 21833 23511
rect 21508 23480 21833 23508
rect 21508 23468 21514 23480
rect 21821 23477 21833 23480
rect 21867 23477 21879 23511
rect 21821 23471 21879 23477
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 23017 23511 23075 23517
rect 23017 23508 23029 23511
rect 22980 23480 23029 23508
rect 22980 23468 22986 23480
rect 23017 23477 23029 23480
rect 23063 23508 23075 23511
rect 25498 23508 25504 23520
rect 23063 23480 25504 23508
rect 23063 23477 23075 23480
rect 23017 23471 23075 23477
rect 25498 23468 25504 23480
rect 25556 23468 25562 23520
rect 37369 23511 37427 23517
rect 37369 23477 37381 23511
rect 37415 23508 37427 23511
rect 37918 23508 37924 23520
rect 37415 23480 37924 23508
rect 37415 23477 37427 23480
rect 37369 23471 37427 23477
rect 37918 23468 37924 23480
rect 37976 23468 37982 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 2038 23264 2044 23316
rect 2096 23304 2102 23316
rect 2593 23307 2651 23313
rect 2593 23304 2605 23307
rect 2096 23276 2605 23304
rect 2096 23264 2102 23276
rect 2593 23273 2605 23276
rect 2639 23273 2651 23307
rect 2593 23267 2651 23273
rect 23017 23307 23075 23313
rect 23017 23273 23029 23307
rect 23063 23304 23075 23307
rect 23290 23304 23296 23316
rect 23063 23276 23296 23304
rect 23063 23273 23075 23276
rect 23017 23267 23075 23273
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 28074 23264 28080 23316
rect 28132 23304 28138 23316
rect 35526 23304 35532 23316
rect 28132 23276 35532 23304
rect 28132 23264 28138 23276
rect 35526 23264 35532 23276
rect 35584 23264 35590 23316
rect 35618 23236 35624 23248
rect 20732 23208 35624 23236
rect 1854 23100 1860 23112
rect 1815 23072 1860 23100
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 6546 23100 6552 23112
rect 2731 23072 6552 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 6546 23060 6552 23072
rect 6604 23060 6610 23112
rect 19426 23060 19432 23112
rect 19484 23100 19490 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19484 23072 19533 23100
rect 19484 23060 19490 23072
rect 19521 23069 19533 23072
rect 19567 23100 19579 23103
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 19567 23072 20637 23100
rect 19567 23069 19579 23072
rect 19521 23063 19579 23069
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 19334 23032 19340 23044
rect 17368 23004 19340 23032
rect 17368 22992 17374 23004
rect 19334 22992 19340 23004
rect 19392 23032 19398 23044
rect 19889 23035 19947 23041
rect 19889 23032 19901 23035
rect 19392 23004 19901 23032
rect 19392 22992 19398 23004
rect 19889 23001 19901 23004
rect 19935 23032 19947 23035
rect 20732 23032 20760 23208
rect 35618 23196 35624 23208
rect 35676 23236 35682 23248
rect 37274 23236 37280 23248
rect 35676 23208 37280 23236
rect 35676 23196 35682 23208
rect 37274 23196 37280 23208
rect 37332 23196 37338 23248
rect 21913 23171 21971 23177
rect 21913 23137 21925 23171
rect 21959 23168 21971 23171
rect 22649 23171 22707 23177
rect 22649 23168 22661 23171
rect 21959 23140 22661 23168
rect 21959 23137 21971 23140
rect 21913 23131 21971 23137
rect 22649 23137 22661 23140
rect 22695 23137 22707 23171
rect 37182 23168 37188 23180
rect 37143 23140 37188 23168
rect 22649 23131 22707 23137
rect 37182 23128 37188 23140
rect 37240 23128 37246 23180
rect 37918 23168 37924 23180
rect 37879 23140 37924 23168
rect 37918 23128 37924 23140
rect 37976 23128 37982 23180
rect 38102 23168 38108 23180
rect 38063 23140 38108 23168
rect 38102 23128 38108 23140
rect 38160 23128 38166 23180
rect 21818 23100 21824 23112
rect 21779 23072 21824 23100
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 22094 23060 22100 23112
rect 22152 23100 22158 23112
rect 23109 23103 23167 23109
rect 23109 23100 23121 23103
rect 22152 23072 23121 23100
rect 22152 23060 22158 23072
rect 23109 23069 23121 23072
rect 23155 23100 23167 23103
rect 24578 23100 24584 23112
rect 23155 23072 24584 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 28074 23060 28080 23112
rect 28132 23100 28138 23112
rect 28169 23103 28227 23109
rect 28169 23100 28181 23103
rect 28132 23072 28181 23100
rect 28132 23060 28138 23072
rect 28169 23069 28181 23072
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 19935 23004 20760 23032
rect 20901 23035 20959 23041
rect 19935 23001 19947 23004
rect 19889 22995 19947 23001
rect 20901 23001 20913 23035
rect 20947 23032 20959 23035
rect 21174 23032 21180 23044
rect 20947 23004 21180 23032
rect 20947 23001 20959 23004
rect 20901 22995 20959 23001
rect 21174 22992 21180 23004
rect 21232 22992 21238 23044
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 20990 22964 20996 22976
rect 1995 22936 20996 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 20990 22924 20996 22936
rect 21048 22924 21054 22976
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22189 22967 22247 22973
rect 22189 22964 22201 22967
rect 22152 22936 22201 22964
rect 22152 22924 22158 22936
rect 22189 22933 22201 22936
rect 22235 22933 22247 22967
rect 22189 22927 22247 22933
rect 28261 22967 28319 22973
rect 28261 22933 28273 22967
rect 28307 22964 28319 22967
rect 28350 22964 28356 22976
rect 28307 22936 28356 22964
rect 28307 22933 28319 22936
rect 28261 22927 28319 22933
rect 28350 22924 28356 22936
rect 28408 22924 28414 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 20714 22760 20720 22772
rect 20627 22732 20720 22760
rect 20714 22720 20720 22732
rect 20772 22760 20778 22772
rect 25590 22760 25596 22772
rect 20772 22732 25596 22760
rect 20772 22720 20778 22732
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 20898 22652 20904 22704
rect 20956 22692 20962 22704
rect 23474 22692 23480 22704
rect 20956 22664 21956 22692
rect 20956 22652 20962 22664
rect 21928 22636 21956 22664
rect 22480 22664 23480 22692
rect 19426 22624 19432 22636
rect 19339 22596 19432 22624
rect 19426 22584 19432 22596
rect 19484 22624 19490 22636
rect 19702 22624 19708 22636
rect 19484 22596 19708 22624
rect 19484 22584 19490 22596
rect 19702 22584 19708 22596
rect 19760 22624 19766 22636
rect 20441 22627 20499 22633
rect 20441 22624 20453 22627
rect 19760 22596 20453 22624
rect 19760 22584 19766 22596
rect 20441 22593 20453 22596
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21140 22596 21833 22624
rect 21140 22584 21146 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22480 22633 22508 22664
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 28350 22692 28356 22704
rect 28311 22664 28356 22692
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21968 22596 22017 22624
rect 21968 22584 21974 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22554 22584 22560 22636
rect 22612 22624 22618 22636
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 22612 22596 22661 22624
rect 22612 22584 22618 22596
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 28166 22624 28172 22636
rect 28127 22596 28172 22624
rect 22649 22587 22707 22593
rect 28166 22584 28172 22596
rect 28224 22584 28230 22636
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22624 37611 22627
rect 37734 22624 37740 22636
rect 37599 22596 37740 22624
rect 37599 22593 37611 22596
rect 37553 22587 37611 22593
rect 37734 22584 37740 22596
rect 37792 22584 37798 22636
rect 19613 22559 19671 22565
rect 19613 22525 19625 22559
rect 19659 22556 19671 22559
rect 20254 22556 20260 22568
rect 19659 22528 20260 22556
rect 19659 22525 19671 22528
rect 19613 22519 19671 22525
rect 20254 22516 20260 22528
rect 20312 22516 20318 22568
rect 30006 22556 30012 22568
rect 29967 22528 30012 22556
rect 30006 22516 30012 22528
rect 30064 22516 30070 22568
rect 22002 22420 22008 22432
rect 21963 22392 22008 22420
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 22462 22380 22468 22432
rect 22520 22420 22526 22432
rect 22557 22423 22615 22429
rect 22557 22420 22569 22423
rect 22520 22392 22569 22420
rect 22520 22380 22526 22392
rect 22557 22389 22569 22392
rect 22603 22389 22615 22423
rect 36538 22420 36544 22432
rect 36499 22392 36544 22420
rect 22557 22383 22615 22389
rect 36538 22380 36544 22392
rect 36596 22380 36602 22432
rect 36630 22380 36636 22432
rect 36688 22420 36694 22432
rect 37645 22423 37703 22429
rect 37645 22420 37657 22423
rect 36688 22392 37657 22420
rect 36688 22380 36694 22392
rect 37645 22389 37657 22392
rect 37691 22389 37703 22423
rect 37645 22383 37703 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 22465 22219 22523 22225
rect 22465 22216 22477 22219
rect 22066 22188 22477 22216
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 22066 22148 22094 22188
rect 22465 22185 22477 22188
rect 22511 22216 22523 22219
rect 23842 22216 23848 22228
rect 22511 22188 23848 22216
rect 22511 22185 22523 22188
rect 22465 22179 22523 22185
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 21876 22120 22094 22148
rect 21876 22108 21882 22120
rect 22557 22083 22615 22089
rect 22557 22049 22569 22083
rect 22603 22080 22615 22083
rect 23474 22080 23480 22092
rect 22603 22052 23480 22080
rect 22603 22049 22615 22052
rect 22557 22043 22615 22049
rect 23474 22040 23480 22052
rect 23532 22080 23538 22092
rect 24026 22080 24032 22092
rect 23532 22052 24032 22080
rect 23532 22040 23538 22052
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 36265 22083 36323 22089
rect 36265 22049 36277 22083
rect 36311 22080 36323 22083
rect 36538 22080 36544 22092
rect 36311 22052 36544 22080
rect 36311 22049 36323 22052
rect 36265 22043 36323 22049
rect 36538 22040 36544 22052
rect 36596 22040 36602 22092
rect 38102 22080 38108 22092
rect 38063 22052 38108 22080
rect 38102 22040 38108 22052
rect 38160 22040 38166 22092
rect 19702 22012 19708 22024
rect 19663 21984 19708 22012
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 20162 22012 20168 22024
rect 20123 21984 20168 22012
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 22002 21972 22008 22024
rect 22060 22021 22066 22024
rect 22060 22015 22096 22021
rect 22084 21981 22096 22015
rect 22060 21975 22096 21981
rect 22060 21972 22066 21975
rect 19426 21944 19432 21956
rect 19387 21916 19432 21944
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 36449 21947 36507 21953
rect 36449 21913 36461 21947
rect 36495 21944 36507 21947
rect 36630 21944 36636 21956
rect 36495 21916 36636 21944
rect 36495 21913 36507 21916
rect 36449 21907 36507 21913
rect 36630 21904 36636 21916
rect 36688 21904 36694 21956
rect 21913 21879 21971 21885
rect 21913 21845 21925 21879
rect 21959 21876 21971 21879
rect 22002 21876 22008 21888
rect 21959 21848 22008 21876
rect 21959 21845 21971 21848
rect 21913 21839 21971 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22186 21876 22192 21888
rect 22143 21848 22192 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22186 21836 22192 21848
rect 22244 21876 22250 21888
rect 23566 21876 23572 21888
rect 22244 21848 23572 21876
rect 22244 21836 22250 21848
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19484 21508 19717 21536
rect 19484 21496 19490 21508
rect 19705 21505 19717 21508
rect 19751 21536 19763 21539
rect 20254 21536 20260 21548
rect 19751 21508 20260 21536
rect 19751 21505 19763 21508
rect 19705 21499 19763 21505
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21536 22063 21539
rect 22186 21536 22192 21548
rect 22051 21508 22192 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21536 23075 21539
rect 23474 21536 23480 21548
rect 23063 21508 23480 21536
rect 23063 21505 23075 21508
rect 23017 21499 23075 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 31754 21496 31760 21548
rect 31812 21536 31818 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 31812 21508 37473 21536
rect 31812 21496 31818 21508
rect 37461 21505 37473 21508
rect 37507 21536 37519 21539
rect 37642 21536 37648 21548
rect 37507 21508 37648 21536
rect 37507 21505 37519 21508
rect 37461 21499 37519 21505
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 21910 21468 21916 21480
rect 21871 21440 21916 21468
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 22925 21471 22983 21477
rect 22925 21468 22937 21471
rect 22388 21440 22937 21468
rect 22388 21409 22416 21440
rect 22925 21437 22937 21440
rect 22971 21437 22983 21471
rect 22925 21431 22983 21437
rect 22373 21403 22431 21409
rect 22373 21369 22385 21403
rect 22419 21369 22431 21403
rect 23382 21400 23388 21412
rect 23343 21372 23388 21400
rect 22373 21363 22431 21369
rect 23382 21360 23388 21372
rect 23440 21360 23446 21412
rect 19794 21332 19800 21344
rect 19755 21304 19800 21332
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 20438 21332 20444 21344
rect 20036 21304 20444 21332
rect 20036 21292 20042 21304
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 36262 21292 36268 21344
rect 36320 21332 36326 21344
rect 36541 21335 36599 21341
rect 36541 21332 36553 21335
rect 36320 21304 36553 21332
rect 36320 21292 36326 21304
rect 36541 21301 36553 21304
rect 36587 21301 36599 21335
rect 36541 21295 36599 21301
rect 36630 21292 36636 21344
rect 36688 21332 36694 21344
rect 37553 21335 37611 21341
rect 37553 21332 37565 21335
rect 36688 21304 37565 21332
rect 36688 21292 36694 21304
rect 37553 21301 37565 21304
rect 37599 21301 37611 21335
rect 37553 21295 37611 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 20346 21020 20352 21072
rect 20404 21060 20410 21072
rect 20404 21032 24624 21060
rect 20404 21020 20410 21032
rect 19981 20995 20039 21001
rect 19981 20961 19993 20995
rect 20027 20992 20039 20995
rect 20162 20992 20168 21004
rect 20027 20964 20168 20992
rect 20027 20961 20039 20964
rect 19981 20955 20039 20961
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 22060 20964 22385 20992
rect 22060 20952 22066 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 22462 20924 22468 20936
rect 22423 20896 22468 20924
rect 22462 20884 22468 20896
rect 22520 20884 22526 20936
rect 24596 20933 24624 21032
rect 36262 20992 36268 21004
rect 36223 20964 36268 20992
rect 36262 20952 36268 20964
rect 36320 20952 36326 21004
rect 36449 20995 36507 21001
rect 36449 20961 36461 20995
rect 36495 20992 36507 20995
rect 36630 20992 36636 21004
rect 36495 20964 36636 20992
rect 36495 20961 36507 20964
rect 36449 20955 36507 20961
rect 36630 20952 36636 20964
rect 36688 20952 36694 21004
rect 38102 20992 38108 21004
rect 38063 20964 38108 20992
rect 38102 20952 38108 20964
rect 38160 20952 38166 21004
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20924 24639 20927
rect 31754 20924 31760 20936
rect 24627 20896 31760 20924
rect 24627 20893 24639 20896
rect 24581 20887 24639 20893
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 20165 20859 20223 20865
rect 20165 20856 20177 20859
rect 19852 20828 20177 20856
rect 19852 20816 19858 20828
rect 20165 20825 20177 20828
rect 20211 20825 20223 20859
rect 20165 20819 20223 20825
rect 21821 20859 21879 20865
rect 21821 20825 21833 20859
rect 21867 20856 21879 20859
rect 34514 20856 34520 20868
rect 21867 20828 34520 20856
rect 21867 20825 21879 20828
rect 21821 20819 21879 20825
rect 34514 20816 34520 20828
rect 34572 20816 34578 20868
rect 22833 20791 22891 20797
rect 22833 20757 22845 20791
rect 22879 20788 22891 20791
rect 23198 20788 23204 20800
rect 22879 20760 23204 20788
rect 22879 20757 22891 20760
rect 22833 20751 22891 20757
rect 23198 20748 23204 20760
rect 23256 20748 23262 20800
rect 24210 20748 24216 20800
rect 24268 20788 24274 20800
rect 24489 20791 24547 20797
rect 24489 20788 24501 20791
rect 24268 20760 24501 20788
rect 24268 20748 24274 20760
rect 24489 20757 24501 20760
rect 24535 20757 24547 20791
rect 24489 20751 24547 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23017 20587 23075 20593
rect 23017 20584 23029 20587
rect 22980 20556 23029 20584
rect 22980 20544 22986 20556
rect 23017 20553 23029 20556
rect 23063 20553 23075 20587
rect 23198 20584 23204 20596
rect 23159 20556 23204 20584
rect 23017 20547 23075 20553
rect 23198 20544 23204 20556
rect 23256 20544 23262 20596
rect 2130 20476 2136 20528
rect 2188 20516 2194 20528
rect 2188 20488 2774 20516
rect 2188 20476 2194 20488
rect 2222 20448 2228 20460
rect 2183 20420 2228 20448
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2746 20448 2774 20488
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 23109 20519 23167 20525
rect 23109 20516 23121 20519
rect 22152 20488 23121 20516
rect 22152 20476 22158 20488
rect 23109 20485 23121 20488
rect 23155 20485 23167 20519
rect 23382 20516 23388 20528
rect 23343 20488 23388 20516
rect 23109 20479 23167 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 24210 20516 24216 20528
rect 24171 20488 24216 20516
rect 24210 20476 24216 20488
rect 24268 20476 24274 20528
rect 25424 20488 26234 20516
rect 2869 20451 2927 20457
rect 2869 20448 2881 20451
rect 2746 20420 2881 20448
rect 2869 20417 2881 20420
rect 2915 20448 2927 20451
rect 21174 20448 21180 20460
rect 2915 20420 21180 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 21174 20408 21180 20420
rect 21232 20448 21238 20460
rect 22002 20448 22008 20460
rect 21232 20420 22008 20448
rect 21232 20408 21238 20420
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 23400 20448 23428 20476
rect 24029 20451 24087 20457
rect 24029 20448 24041 20451
rect 23400 20420 24041 20448
rect 24029 20417 24041 20420
rect 24075 20417 24087 20451
rect 24029 20411 24087 20417
rect 18598 20340 18604 20392
rect 18656 20380 18662 20392
rect 25424 20380 25452 20488
rect 26206 20448 26234 20488
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 26206 20420 37473 20448
rect 37461 20417 37473 20420
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 25866 20380 25872 20392
rect 18656 20352 25452 20380
rect 25827 20352 25872 20380
rect 18656 20340 18662 20352
rect 25866 20340 25872 20352
rect 25924 20340 25930 20392
rect 21358 20272 21364 20324
rect 21416 20312 21422 20324
rect 22833 20315 22891 20321
rect 22833 20312 22845 20315
rect 21416 20284 22845 20312
rect 21416 20272 21422 20284
rect 22833 20281 22845 20284
rect 22879 20281 22891 20315
rect 22833 20275 22891 20281
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 1670 20244 1676 20256
rect 1627 20216 1676 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 1670 20204 1676 20216
rect 1728 20204 1734 20256
rect 2130 20244 2136 20256
rect 2091 20216 2136 20244
rect 2130 20204 2136 20216
rect 2188 20204 2194 20256
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 22097 20247 22155 20253
rect 2832 20216 2877 20244
rect 2832 20204 2838 20216
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22186 20244 22192 20256
rect 22143 20216 22192 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 37553 20247 37611 20253
rect 37553 20213 37565 20247
rect 37599 20244 37611 20247
rect 37918 20244 37924 20256
rect 37599 20216 37924 20244
rect 37599 20213 37611 20216
rect 37553 20207 37611 20213
rect 37918 20204 37924 20216
rect 37976 20204 37982 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2130 19972 2136 19984
rect 1596 19944 2136 19972
rect 1596 19913 1624 19944
rect 2130 19932 2136 19944
rect 2188 19932 2194 19984
rect 22094 19972 22100 19984
rect 22020 19944 22100 19972
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19873 1639 19907
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1581 19867 1639 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 22020 19913 22048 19944
rect 22094 19932 22100 19944
rect 22152 19932 22158 19984
rect 22005 19907 22063 19913
rect 22005 19873 22017 19907
rect 22051 19873 22063 19907
rect 22186 19904 22192 19916
rect 22147 19876 22192 19904
rect 22005 19867 22063 19873
rect 22186 19864 22192 19876
rect 22244 19864 22250 19916
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 23256 19876 24409 19904
rect 23256 19864 23262 19876
rect 24397 19873 24409 19876
rect 24443 19873 24455 19907
rect 37182 19904 37188 19916
rect 37143 19876 37188 19904
rect 24397 19867 24455 19873
rect 37182 19864 37188 19876
rect 37240 19864 37246 19916
rect 37918 19904 37924 19916
rect 37879 19876 37924 19904
rect 37918 19864 37924 19876
rect 37976 19864 37982 19916
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 21358 19836 21364 19848
rect 21319 19808 21364 19836
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 31754 19836 31760 19848
rect 31715 19808 31760 19836
rect 31754 19796 31760 19808
rect 31812 19796 31818 19848
rect 38102 19796 38108 19848
rect 38160 19836 38166 19848
rect 38160 19808 38205 19836
rect 38160 19796 38166 19808
rect 23842 19768 23848 19780
rect 23803 19740 23848 19768
rect 23842 19728 23848 19740
rect 23900 19728 23906 19780
rect 24578 19768 24584 19780
rect 24539 19740 24584 19768
rect 24578 19728 24584 19740
rect 24636 19728 24642 19780
rect 26237 19771 26295 19777
rect 26237 19737 26249 19771
rect 26283 19768 26295 19771
rect 35618 19768 35624 19780
rect 26283 19740 35624 19768
rect 26283 19737 26295 19740
rect 26237 19731 26295 19737
rect 35618 19728 35624 19740
rect 35676 19728 35682 19780
rect 21545 19703 21603 19709
rect 21545 19669 21557 19703
rect 21591 19700 21603 19703
rect 22094 19700 22100 19712
rect 21591 19672 22100 19700
rect 21591 19669 21603 19672
rect 21545 19663 21603 19669
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 31849 19703 31907 19709
rect 31849 19669 31861 19703
rect 31895 19700 31907 19703
rect 32306 19700 32312 19712
rect 31895 19672 32312 19700
rect 31895 19669 31907 19672
rect 31849 19663 31907 19669
rect 32306 19660 32312 19672
rect 32364 19660 32370 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 24489 19499 24547 19505
rect 24489 19465 24501 19499
rect 24535 19496 24547 19499
rect 24578 19496 24584 19508
rect 24535 19468 24584 19496
rect 24535 19465 24547 19468
rect 24489 19459 24547 19465
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 1857 19431 1915 19437
rect 1857 19397 1869 19431
rect 1903 19428 1915 19431
rect 2774 19428 2780 19440
rect 1903 19400 2780 19428
rect 1903 19397 1915 19400
rect 1857 19391 1915 19397
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 32306 19428 32312 19440
rect 22060 19400 24440 19428
rect 32267 19400 32312 19428
rect 22060 19388 22066 19400
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 22094 19360 22100 19372
rect 22055 19332 22100 19360
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 23934 19360 23940 19372
rect 23895 19332 23940 19360
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24412 19369 24440 19400
rect 32306 19388 32312 19400
rect 32364 19388 32370 19440
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19329 24455 19363
rect 24397 19323 24455 19329
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19360 37887 19363
rect 38102 19360 38108 19372
rect 37875 19332 38108 19360
rect 37875 19329 37887 19332
rect 37829 19323 37887 19329
rect 38102 19320 38108 19332
rect 38160 19320 38166 19372
rect 2130 19292 2136 19304
rect 2091 19264 2136 19292
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 22278 19292 22284 19304
rect 22239 19264 22284 19292
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 31573 19295 31631 19301
rect 31573 19261 31585 19295
rect 31619 19292 31631 19295
rect 32125 19295 32183 19301
rect 32125 19292 32137 19295
rect 31619 19264 32137 19292
rect 31619 19261 31631 19264
rect 31573 19255 31631 19261
rect 32125 19261 32137 19264
rect 32171 19261 32183 19295
rect 32125 19255 32183 19261
rect 32585 19295 32643 19301
rect 32585 19261 32597 19295
rect 32631 19261 32643 19295
rect 32585 19255 32643 19261
rect 31754 19184 31760 19236
rect 31812 19224 31818 19236
rect 32600 19224 32628 19255
rect 31812 19196 32628 19224
rect 31812 19184 31818 19196
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 1673 18955 1731 18961
rect 1673 18952 1685 18955
rect 1452 18924 1685 18952
rect 1452 18912 1458 18924
rect 1673 18921 1685 18924
rect 1719 18921 1731 18955
rect 1673 18915 1731 18921
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 21821 18819 21879 18825
rect 21821 18816 21833 18819
rect 12492 18788 21833 18816
rect 12492 18776 12498 18788
rect 21821 18785 21833 18788
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 20809 18683 20867 18689
rect 20809 18649 20821 18683
rect 20855 18680 20867 18683
rect 21545 18683 21603 18689
rect 21545 18680 21557 18683
rect 20855 18652 21557 18680
rect 20855 18649 20867 18652
rect 20809 18643 20867 18649
rect 21545 18649 21557 18652
rect 21591 18649 21603 18683
rect 21545 18643 21603 18649
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 22278 18408 22284 18420
rect 22239 18380 22284 18408
rect 22278 18368 22284 18380
rect 22336 18368 22342 18420
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 20772 18244 22201 18272
rect 20772 18232 20778 18244
rect 22189 18241 22201 18244
rect 22235 18272 22247 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 22235 18244 26985 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 27065 18071 27123 18077
rect 27065 18037 27077 18071
rect 27111 18068 27123 18071
rect 27246 18068 27252 18080
rect 27111 18040 27252 18068
rect 27111 18037 27123 18040
rect 27065 18031 27123 18037
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 27614 18068 27620 18080
rect 27575 18040 27620 18068
rect 27614 18028 27620 18040
rect 27672 18028 27678 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 27614 17796 27620 17808
rect 27080 17768 27620 17796
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1578 17728 1584 17740
rect 1443 17700 1584 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 27080 17737 27108 17768
rect 27614 17756 27620 17768
rect 27672 17756 27678 17808
rect 27065 17731 27123 17737
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 27065 17697 27077 17731
rect 27111 17697 27123 17731
rect 27246 17728 27252 17740
rect 27207 17700 27252 17728
rect 27065 17691 27123 17697
rect 27246 17688 27252 17700
rect 27304 17688 27310 17740
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 1946 17592 1952 17604
rect 1627 17564 1952 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 28902 17592 28908 17604
rect 28863 17564 28908 17592
rect 28902 17552 28908 17564
rect 28960 17552 28966 17604
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 28353 17255 28411 17261
rect 28353 17221 28365 17255
rect 28399 17252 28411 17255
rect 29089 17255 29147 17261
rect 29089 17252 29101 17255
rect 28399 17224 29101 17252
rect 28399 17221 28411 17224
rect 28353 17215 28411 17221
rect 29089 17221 29101 17224
rect 29135 17221 29147 17255
rect 29089 17215 29147 17221
rect 2038 17184 2044 17196
rect 1951 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17184 2102 17196
rect 9122 17184 9128 17196
rect 2096 17156 9128 17184
rect 2096 17144 2102 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 28261 17187 28319 17193
rect 28261 17184 28273 17187
rect 20680 17156 28273 17184
rect 20680 17144 20686 17156
rect 28261 17153 28273 17156
rect 28307 17153 28319 17187
rect 28261 17147 28319 17153
rect 28905 17119 28963 17125
rect 28905 17085 28917 17119
rect 28951 17116 28963 17119
rect 29546 17116 29552 17128
rect 28951 17088 29552 17116
rect 28951 17085 28963 17088
rect 28905 17079 28963 17085
rect 29546 17076 29552 17088
rect 29604 17076 29610 17128
rect 30745 17119 30803 17125
rect 30745 17085 30757 17119
rect 30791 17116 30803 17119
rect 34514 17116 34520 17128
rect 30791 17088 34520 17116
rect 30791 17085 30803 17088
rect 30745 17079 30803 17085
rect 34514 17076 34520 17088
rect 34572 17076 34578 17128
rect 3602 16980 3608 16992
rect 3563 16952 3608 16980
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 37829 16983 37887 16989
rect 37829 16949 37841 16983
rect 37875 16980 37887 16983
rect 38102 16980 38108 16992
rect 37875 16952 38108 16980
rect 37875 16949 37887 16952
rect 37829 16943 37887 16949
rect 38102 16940 38108 16952
rect 38160 16940 38166 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 29546 16776 29552 16788
rect 29507 16748 29552 16776
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 20622 16708 20628 16720
rect 9508 16680 20628 16708
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 3418 16572 3424 16584
rect 2823 16544 3424 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 2148 16504 2176 16535
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16572 3847 16575
rect 9508 16572 9536 16680
rect 20622 16668 20628 16680
rect 20680 16668 20686 16720
rect 19334 16640 19340 16652
rect 3835 16544 9536 16572
rect 9646 16612 19340 16640
rect 3835 16541 3847 16544
rect 3789 16535 3847 16541
rect 9646 16504 9674 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 37642 16640 37648 16652
rect 37603 16612 37648 16640
rect 37642 16600 37648 16612
rect 37700 16600 37706 16652
rect 38102 16640 38108 16652
rect 38063 16612 38108 16640
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 2148 16476 9674 16504
rect 37550 16464 37556 16516
rect 37608 16504 37614 16516
rect 37921 16507 37979 16513
rect 37921 16504 37933 16507
rect 37608 16476 37933 16504
rect 37608 16464 37614 16476
rect 37921 16473 37933 16476
rect 37967 16473 37979 16507
rect 37921 16467 37979 16473
rect 2041 16439 2099 16445
rect 2041 16405 2053 16439
rect 2087 16436 2099 16439
rect 3234 16436 3240 16448
rect 2087 16408 3240 16436
rect 2087 16405 2099 16408
rect 2041 16399 2099 16405
rect 3234 16396 3240 16408
rect 3292 16396 3298 16448
rect 3881 16439 3939 16445
rect 3881 16405 3893 16439
rect 3927 16436 3939 16439
rect 4062 16436 4068 16448
rect 3927 16408 4068 16436
rect 3927 16405 3939 16408
rect 3881 16399 3939 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 37550 16232 37556 16244
rect 37511 16204 37556 16232
rect 37550 16192 37556 16204
rect 37608 16192 37614 16244
rect 3234 16164 3240 16176
rect 3195 16136 3240 16164
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 4062 16164 4068 16176
rect 4023 16136 4068 16164
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3476 16068 3521 16096
rect 3476 16056 3482 16068
rect 3602 16056 3608 16108
rect 3660 16096 3666 16108
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3660 16068 3893 16096
rect 3660 16056 3666 16068
rect 3881 16065 3893 16068
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 19058 16056 19064 16108
rect 19116 16096 19122 16108
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 19116 16068 37473 16096
rect 19116 16056 19122 16068
rect 37461 16065 37473 16068
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 3436 16000 4353 16028
rect 3436 15972 3464 16000
rect 4341 15997 4353 16000
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 3418 15920 3424 15972
rect 3476 15920 3482 15972
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 4430 15552 4436 15564
rect 2823 15524 4436 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 19058 15552 19064 15564
rect 12406 15524 19064 15552
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15484 4031 15487
rect 12406 15484 12434 15524
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 4019 15456 12434 15484
rect 37829 15487 37887 15493
rect 4019 15453 4031 15456
rect 3973 15447 4031 15453
rect 37829 15453 37841 15487
rect 37875 15484 37887 15487
rect 38102 15484 38108 15496
rect 37875 15456 38108 15484
rect 37875 15453 37887 15456
rect 37829 15447 37887 15453
rect 38102 15444 38108 15456
rect 38160 15444 38166 15496
rect 21818 15416 21824 15428
rect 1596 15388 21824 15416
rect 1596 15357 1624 15388
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4246 15348 4252 15360
rect 3927 15320 4252 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 4246 15076 4252 15088
rect 4207 15048 4252 15076
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2130 15008 2136 15020
rect 2087 14980 2136 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 4430 14968 4436 15020
rect 4488 15008 4494 15020
rect 4488 14980 4533 15008
rect 4488 14968 4494 14980
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 18012 14980 37473 15008
rect 18012 14968 18018 14980
rect 37461 14977 37473 14980
rect 37507 15008 37519 15011
rect 37642 15008 37648 15020
rect 37507 14980 37648 15008
rect 37507 14977 37519 14980
rect 37461 14971 37519 14977
rect 37642 14968 37648 14980
rect 37700 14968 37706 15020
rect 2866 14940 2872 14952
rect 2827 14912 2872 14940
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 1949 14807 2007 14813
rect 1949 14773 1961 14807
rect 1995 14804 2007 14807
rect 3050 14804 3056 14816
rect 1995 14776 3056 14804
rect 1995 14773 2007 14776
rect 1949 14767 2007 14773
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 19794 14804 19800 14816
rect 19755 14776 19800 14804
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 37553 14807 37611 14813
rect 37553 14773 37565 14807
rect 37599 14804 37611 14807
rect 37918 14804 37924 14816
rect 37599 14776 37924 14804
rect 37599 14773 37611 14776
rect 37553 14767 37611 14773
rect 37918 14764 37924 14776
rect 37976 14764 37982 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 19794 14464 19800 14476
rect 19755 14436 19800 14464
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 37182 14464 37188 14476
rect 37143 14436 37188 14464
rect 37182 14424 37188 14436
rect 37240 14424 37246 14476
rect 37918 14464 37924 14476
rect 37879 14436 37924 14464
rect 37918 14424 37924 14436
rect 37976 14424 37982 14476
rect 38102 14464 38108 14476
rect 38063 14436 38108 14464
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3283 14368 3801 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19981 14331 20039 14337
rect 19981 14328 19993 14331
rect 19484 14300 19993 14328
rect 19484 14288 19490 14300
rect 19981 14297 19993 14300
rect 20027 14297 20039 14331
rect 19981 14291 20039 14297
rect 21637 14331 21695 14337
rect 21637 14297 21649 14331
rect 21683 14328 21695 14331
rect 34514 14328 34520 14340
rect 21683 14300 34520 14328
rect 21683 14297 21695 14300
rect 21637 14291 21695 14297
rect 34514 14288 34520 14300
rect 34572 14288 34578 14340
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 18690 13880 18696 13932
rect 18748 13920 18754 13932
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 18748 13892 19349 13920
rect 18748 13880 18754 13892
rect 19337 13889 19349 13892
rect 19383 13920 19395 13923
rect 19426 13920 19432 13932
rect 19383 13892 19432 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 3510 13852 3516 13864
rect 3471 13824 3516 13852
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3694 13852 3700 13864
rect 3655 13824 3700 13852
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 37826 13716 37832 13728
rect 37787 13688 37832 13716
rect 37826 13676 37832 13688
rect 37884 13676 37890 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2593 13515 2651 13521
rect 2593 13481 2605 13515
rect 2639 13512 2651 13515
rect 3510 13512 3516 13524
rect 2639 13484 3516 13512
rect 2639 13481 2651 13484
rect 2593 13475 2651 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 37182 13376 37188 13388
rect 37143 13348 37188 13376
rect 37182 13336 37188 13348
rect 37240 13336 37246 13388
rect 37826 13336 37832 13388
rect 37884 13376 37890 13388
rect 38105 13379 38163 13385
rect 38105 13376 38117 13379
rect 37884 13348 38117 13376
rect 37884 13336 37890 13348
rect 38105 13345 38117 13348
rect 38151 13345 38163 13379
rect 38105 13339 38163 13345
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1452 13280 1593 13308
rect 1452 13268 1458 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13308 2743 13311
rect 2731 13280 4016 13308
rect 2731 13277 2743 13280
rect 2685 13271 2743 13277
rect 3988 13184 4016 13280
rect 37550 13200 37556 13252
rect 37608 13240 37614 13252
rect 37921 13243 37979 13249
rect 37921 13240 37933 13243
rect 37608 13212 37933 13240
rect 37608 13200 37614 13212
rect 37921 13209 37933 13212
rect 37967 13209 37979 13243
rect 37921 13203 37979 13209
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 19426 13172 19432 13184
rect 4028 13144 19432 13172
rect 4028 13132 4034 13144
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 37550 12968 37556 12980
rect 37511 12940 37556 12968
rect 37550 12928 37556 12940
rect 37608 12928 37614 12980
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2222 12832 2228 12844
rect 2087 12804 2228 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 3694 12832 3700 12844
rect 2731 12804 3700 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 20254 12832 20260 12844
rect 12406 12804 20260 12832
rect 2240 12764 2268 12792
rect 12406 12764 12434 12804
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 37458 12832 37464 12844
rect 37371 12804 37464 12832
rect 37458 12792 37464 12804
rect 37516 12832 37522 12844
rect 37734 12832 37740 12844
rect 37516 12804 37740 12832
rect 37516 12792 37522 12804
rect 37734 12792 37740 12804
rect 37792 12792 37798 12844
rect 2240 12736 12434 12764
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1636 12600 1961 12628
rect 1636 12588 1642 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 1949 12591 2007 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 1578 12288 1584 12300
rect 1539 12260 1584 12288
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 2774 12288 2780 12300
rect 2735 12260 2780 12288
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 37182 12288 37188 12300
rect 37143 12260 37188 12288
rect 37182 12248 37188 12260
rect 37240 12248 37246 12300
rect 35802 12180 35808 12232
rect 35860 12220 35866 12232
rect 36265 12223 36323 12229
rect 36265 12220 36277 12223
rect 35860 12192 36277 12220
rect 35860 12180 35866 12192
rect 36265 12189 36277 12192
rect 36311 12189 36323 12223
rect 36265 12183 36323 12189
rect 36449 12155 36507 12161
rect 36449 12121 36461 12155
rect 36495 12152 36507 12155
rect 37274 12152 37280 12164
rect 36495 12124 37280 12152
rect 36495 12121 36507 12124
rect 36449 12115 36507 12121
rect 37274 12112 37280 12124
rect 37332 12112 37338 12164
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 37826 11744 37832 11756
rect 37599 11716 37832 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 37826 11704 37832 11716
rect 37884 11704 37890 11756
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2038 11676 2044 11688
rect 1903 11648 2044 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 36262 11500 36268 11552
rect 36320 11540 36326 11552
rect 36541 11543 36599 11549
rect 36541 11540 36553 11543
rect 36320 11512 36553 11540
rect 36320 11500 36326 11512
rect 36541 11509 36553 11512
rect 36587 11509 36599 11543
rect 37642 11540 37648 11552
rect 37603 11512 37648 11540
rect 36541 11503 36599 11509
rect 37642 11500 37648 11512
rect 37700 11500 37706 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 35802 11336 35808 11348
rect 35763 11308 35808 11336
rect 35802 11296 35808 11308
rect 35860 11296 35866 11348
rect 36262 11200 36268 11212
rect 36223 11172 36268 11200
rect 36262 11160 36268 11172
rect 36320 11160 36326 11212
rect 36449 11203 36507 11209
rect 36449 11169 36461 11203
rect 36495 11200 36507 11203
rect 37642 11200 37648 11212
rect 36495 11172 37648 11200
rect 36495 11169 36507 11172
rect 36449 11163 36507 11169
rect 37642 11160 37648 11172
rect 37700 11160 37706 11212
rect 38102 11200 38108 11212
rect 38063 11172 38108 11200
rect 38102 11160 38108 11172
rect 38160 11160 38166 11212
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2682 11132 2688 11144
rect 2179 11104 2688 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2682 11092 2688 11104
rect 2740 11132 2746 11144
rect 18138 11132 18144 11144
rect 2740 11104 18144 11132
rect 2740 11092 2746 11104
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 18564 11104 19717 11132
rect 18564 11092 18570 11104
rect 19705 11101 19717 11104
rect 19751 11132 19763 11135
rect 20162 11132 20168 11144
rect 19751 11104 20168 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 20162 11092 20168 11104
rect 20220 11092 20226 11144
rect 20254 11064 20260 11076
rect 20167 11036 20260 11064
rect 20254 11024 20260 11036
rect 20312 11064 20318 11076
rect 37826 11064 37832 11076
rect 20312 11036 37832 11064
rect 20312 11024 20318 11036
rect 37826 11024 37832 11036
rect 37884 11024 37890 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 37274 10752 37280 10804
rect 37332 10792 37338 10804
rect 37553 10795 37611 10801
rect 37553 10792 37565 10795
rect 37332 10764 37565 10792
rect 37332 10752 37338 10764
rect 37553 10761 37565 10764
rect 37599 10761 37611 10795
rect 37553 10755 37611 10761
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6546 10616 6552 10628
rect 6604 10656 6610 10668
rect 20254 10656 20260 10668
rect 6604 10628 20260 10656
rect 6604 10616 6610 10628
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 37461 10659 37519 10665
rect 37461 10625 37473 10659
rect 37507 10656 37519 10659
rect 37826 10656 37832 10668
rect 37507 10628 37832 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 37826 10616 37832 10628
rect 37884 10616 37890 10668
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6144 10424 6469 10452
rect 6144 10412 6150 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 36262 10412 36268 10464
rect 36320 10452 36326 10464
rect 36541 10455 36599 10461
rect 36541 10452 36553 10455
rect 36320 10424 36553 10452
rect 36320 10412 36326 10424
rect 36541 10421 36553 10424
rect 36587 10421 36599 10455
rect 36541 10415 36599 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6328 10084 6377 10112
rect 6328 10072 6334 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 36262 10112 36268 10124
rect 36223 10084 36268 10112
rect 6365 10075 6423 10081
rect 36262 10072 36268 10084
rect 36320 10072 36326 10124
rect 38102 10112 38108 10124
rect 38063 10084 38108 10112
rect 38102 10072 38108 10084
rect 38160 10072 38166 10124
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5491 10016 5917 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 36446 9976 36452 9988
rect 36407 9948 36452 9976
rect 36446 9936 36452 9948
rect 36504 9936 36510 9988
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 36446 9664 36452 9716
rect 36504 9704 36510 9716
rect 36633 9707 36691 9713
rect 36633 9704 36645 9707
rect 36504 9676 36645 9704
rect 36504 9664 36510 9676
rect 36633 9673 36645 9676
rect 36679 9673 36691 9707
rect 36633 9667 36691 9673
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 36725 9571 36783 9577
rect 36725 9568 36737 9571
rect 18472 9540 36737 9568
rect 18472 9528 18478 9540
rect 36725 9537 36737 9540
rect 36771 9537 36783 9571
rect 37366 9568 37372 9580
rect 37327 9540 37372 9568
rect 36725 9531 36783 9537
rect 37366 9528 37372 9540
rect 37424 9528 37430 9580
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1452 9336 1593 9364
rect 1452 9324 1458 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 37461 9367 37519 9373
rect 37461 9333 37473 9367
rect 37507 9364 37519 9367
rect 37918 9364 37924 9376
rect 37507 9336 37924 9364
rect 37507 9333 37519 9336
rect 37461 9327 37519 9333
rect 37918 9324 37924 9336
rect 37976 9324 37982 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 37182 9024 37188 9036
rect 37143 8996 37188 9024
rect 37182 8984 37188 8996
rect 37240 8984 37246 9036
rect 37918 9024 37924 9036
rect 37879 8996 37924 9024
rect 37918 8984 37924 8996
rect 37976 8984 37982 9036
rect 38102 8916 38108 8968
rect 38160 8956 38166 8968
rect 38160 8928 38205 8956
rect 38160 8916 38166 8928
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 1946 8888 1952 8900
rect 1627 8860 1952 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 1946 8848 1952 8860
rect 2004 8848 2010 8900
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2130 8480 2136 8492
rect 2087 8452 2136 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2682 8480 2688 8492
rect 2643 8452 2688 8480
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 19334 8440 19340 8492
rect 19392 8480 19398 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19392 8452 19993 8480
rect 19392 8440 19398 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8480 37887 8483
rect 38102 8480 38108 8492
rect 37875 8452 38108 8480
rect 37875 8449 37887 8452
rect 37829 8443 37887 8449
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 4212 8384 7941 8412
rect 4212 8372 4218 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 9582 8412 9588 8424
rect 9543 8384 9588 8412
rect 7929 8375 7987 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 3050 8344 3056 8356
rect 2639 8316 3056 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 9784 8344 9812 8375
rect 8352 8316 9812 8344
rect 8352 8304 8358 8316
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3234 8276 3240 8288
rect 3191 8248 3240 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 20073 8279 20131 8285
rect 20073 8245 20085 8279
rect 20119 8276 20131 8279
rect 20622 8276 20628 8288
rect 20119 8248 20628 8276
rect 20119 8245 20131 8248
rect 20073 8239 20131 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8294 8072 8300 8084
rect 8159 8044 8300 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 9582 8072 9588 8084
rect 9079 8044 9588 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 3050 7936 3056 7948
rect 3011 7908 3056 7936
rect 3050 7896 3056 7908
rect 3108 7896 3114 7948
rect 3234 7936 3240 7948
rect 3195 7908 3240 7936
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 20622 7936 20628 7948
rect 20583 7908 20628 7936
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 22002 7936 22008 7948
rect 21963 7908 22008 7936
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 9122 7868 9128 7880
rect 9035 7840 9128 7868
rect 9122 7828 9128 7840
rect 9180 7868 9186 7880
rect 18598 7868 18604 7880
rect 9180 7840 18604 7868
rect 9180 7828 9186 7840
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 1394 7800 1400 7812
rect 1355 7772 1400 7800
rect 1394 7760 1400 7772
rect 1452 7760 1458 7812
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20496 7364 20545 7392
rect 20496 7352 20502 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9398 7188 9404 7200
rect 9263 7160 9404 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 9398 6848 9404 6860
rect 9359 6820 9404 6848
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9232 6712 9260 6743
rect 9766 6712 9772 6724
rect 9232 6684 9772 6712
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 1946 6236 1952 6248
rect 1811 6208 1952 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2038 6196 2044 6248
rect 2096 6236 2102 6248
rect 2096 6208 2141 6236
rect 2096 6196 2102 6208
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2130 5692 2136 5704
rect 2087 5664 2136 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2130 5652 2136 5664
rect 2188 5692 2194 5704
rect 2406 5692 2412 5704
rect 2188 5664 2412 5692
rect 2188 5652 2194 5664
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 23934 5352 23940 5364
rect 3384 5324 23940 5352
rect 3384 5312 3390 5324
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10468 4984 10517 5012
rect 10468 4972 10474 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 10505 4975 10563 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 37829 5015 37887 5021
rect 37829 4981 37841 5015
rect 37875 5012 37887 5015
rect 38102 5012 38108 5024
rect 37875 4984 38108 5012
rect 37875 4981 37887 4984
rect 37829 4975 37887 4981
rect 38102 4972 38108 4984
rect 38160 4972 38166 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 9732 4712 11100 4740
rect 9732 4700 9738 4712
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 3234 4672 3240 4684
rect 1811 4644 3240 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 10410 4672 10416 4684
rect 10371 4644 10416 4672
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 11072 4681 11100 4712
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4641 11115 4675
rect 37182 4672 37188 4684
rect 11057 4635 11115 4641
rect 18616 4644 20300 4672
rect 37143 4644 37188 4672
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 2961 4607 3019 4613
rect 2961 4604 2973 4607
rect 2924 4576 2973 4604
rect 2924 4564 2930 4576
rect 2961 4573 2973 4576
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4604 17923 4607
rect 18506 4604 18512 4616
rect 17911 4576 18512 4604
rect 17911 4573 17923 4576
rect 17865 4567 17923 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18616 4613 18644 4644
rect 20272 4616 20300 4644
rect 37182 4632 37188 4644
rect 37240 4632 37246 4684
rect 38102 4672 38108 4684
rect 38063 4644 38108 4672
rect 38102 4632 38108 4644
rect 38160 4632 38166 4684
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4573 18659 4607
rect 19426 4604 19432 4616
rect 19387 4576 19432 4604
rect 18601 4567 18659 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20312 4576 20729 4604
rect 20312 4564 20318 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20717 4567 20775 4573
rect 10594 4536 10600 4548
rect 10555 4508 10600 4536
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 37918 4536 37924 4548
rect 37879 4508 37924 4536
rect 37918 4496 37924 4508
rect 37976 4496 37982 4548
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18509 4471 18567 4477
rect 18509 4468 18521 4471
rect 18012 4440 18521 4468
rect 18012 4428 18018 4440
rect 18509 4437 18521 4440
rect 18555 4437 18567 4471
rect 20806 4468 20812 4480
rect 20767 4440 20812 4468
rect 18509 4431 18567 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 10505 4267 10563 4273
rect 10505 4233 10517 4267
rect 10551 4264 10563 4267
rect 10594 4264 10600 4276
rect 10551 4236 10600 4264
rect 10551 4233 10563 4236
rect 10505 4227 10563 4233
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 37553 4267 37611 4273
rect 37553 4233 37565 4267
rect 37599 4264 37611 4267
rect 37918 4264 37924 4276
rect 37599 4236 37924 4264
rect 37599 4233 37611 4236
rect 37553 4227 37611 4233
rect 37918 4224 37924 4236
rect 37976 4224 37982 4276
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 17954 4196 17960 4208
rect 3568 4168 17632 4196
rect 17915 4168 17960 4196
rect 3568 4156 3574 4168
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 10410 4128 10416 4140
rect 9999 4100 10416 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3878 4060 3884 4072
rect 3099 4032 3884 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4029 4031 4063
rect 17604 4060 17632 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 36280 4168 36492 4196
rect 17770 4128 17776 4140
rect 17731 4100 17776 4128
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 20622 4128 20628 4140
rect 20583 4100 20628 4128
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 31846 4128 31852 4140
rect 22612 4100 31852 4128
rect 22612 4088 22618 4100
rect 31846 4088 31852 4100
rect 31904 4088 31910 4140
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 36280 4128 36308 4168
rect 35023 4100 36308 4128
rect 36357 4131 36415 4137
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 36357 4097 36369 4131
rect 36403 4097 36415 4131
rect 36464 4128 36492 4168
rect 37274 4128 37280 4140
rect 36464 4100 37280 4128
rect 36357 4091 36415 4097
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 17604 4032 18245 4060
rect 3973 4023 4031 4029
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 34514 4060 34520 4072
rect 18233 4023 18291 4029
rect 26206 4032 34520 4060
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 3988 3992 4016 4023
rect 3384 3964 4016 3992
rect 3384 3952 3390 3964
rect 23658 3952 23664 4004
rect 23716 3992 23722 4004
rect 26206 3992 26234 4032
rect 34514 4020 34520 4032
rect 34572 4020 34578 4072
rect 36372 4060 36400 4091
rect 37274 4088 37280 4100
rect 37332 4128 37338 4140
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 37332 4100 37473 4128
rect 37332 4088 37338 4100
rect 37461 4097 37473 4100
rect 37507 4097 37519 4131
rect 37461 4091 37519 4097
rect 37734 4060 37740 4072
rect 36372 4032 37740 4060
rect 37734 4020 37740 4032
rect 37792 4020 37798 4072
rect 35710 3992 35716 4004
rect 23716 3964 26234 3992
rect 31036 3964 35716 3992
rect 23716 3952 23722 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1673 3927 1731 3933
rect 1673 3924 1685 3927
rect 1452 3896 1685 3924
rect 1452 3884 1458 3896
rect 1673 3893 1685 3896
rect 1719 3893 1731 3927
rect 1673 3887 1731 3893
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 6454 3924 6460 3936
rect 5399 3896 6460 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9364 3896 9873 3924
rect 9364 3884 9370 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 9861 3887 9919 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 21818 3924 21824 3936
rect 21779 3896 21824 3924
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 31036 3924 31064 3964
rect 35710 3952 35716 3964
rect 35768 3952 35774 4004
rect 32306 3924 32312 3936
rect 22336 3896 31064 3924
rect 32267 3896 32312 3924
rect 22336 3884 22342 3896
rect 32306 3884 32312 3896
rect 32364 3884 32370 3936
rect 32582 3884 32588 3936
rect 32640 3924 32646 3936
rect 32953 3927 33011 3933
rect 32953 3924 32965 3927
rect 32640 3896 32965 3924
rect 32640 3884 32646 3896
rect 32953 3893 32965 3896
rect 32999 3893 33011 3927
rect 32953 3887 33011 3893
rect 34057 3927 34115 3933
rect 34057 3893 34069 3927
rect 34103 3924 34115 3927
rect 34698 3924 34704 3936
rect 34103 3896 34704 3924
rect 34103 3893 34115 3896
rect 34057 3887 34115 3893
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 35069 3927 35127 3933
rect 35069 3893 35081 3927
rect 35115 3924 35127 3927
rect 35342 3924 35348 3936
rect 35115 3896 35348 3924
rect 35115 3893 35127 3896
rect 35069 3887 35127 3893
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 35618 3924 35624 3936
rect 35579 3896 35624 3924
rect 35618 3884 35624 3896
rect 35676 3884 35682 3936
rect 36449 3927 36507 3933
rect 36449 3893 36461 3927
rect 36495 3924 36507 3927
rect 37826 3924 37832 3936
rect 36495 3896 37832 3924
rect 36495 3893 36507 3896
rect 36449 3887 36507 3893
rect 37826 3884 37832 3896
rect 37884 3884 37890 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 19981 3723 20039 3729
rect 6886 3692 14504 3720
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 6886 3652 6914 3692
rect 716 3624 6914 3652
rect 8956 3624 9628 3652
rect 716 3612 722 3624
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 2866 3584 2872 3596
rect 2823 3556 2872 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3234 3584 3240 3596
rect 3195 3556 3240 3584
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8662 3516 8668 3528
rect 8159 3488 8668 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 3053 3451 3111 3457
rect 3053 3448 3065 3451
rect 2740 3420 3065 3448
rect 2740 3408 2746 3420
rect 3053 3417 3065 3420
rect 3099 3417 3111 3451
rect 4614 3448 4620 3460
rect 4575 3420 4620 3448
rect 3053 3411 3111 3417
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6273 3451 6331 3457
rect 6273 3448 6285 3451
rect 5776 3420 6285 3448
rect 5776 3408 5782 3420
rect 6273 3417 6285 3420
rect 6319 3417 6331 3451
rect 6273 3411 6331 3417
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 8956 3380 8984 3624
rect 9122 3584 9128 3596
rect 9083 3556 9128 3584
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9600 3593 9628 3624
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14332 3488 14381 3516
rect 14332 3476 14338 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 14476 3516 14504 3692
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20162 3720 20168 3732
rect 20027 3692 20168 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20162 3680 20168 3692
rect 20220 3720 20226 3732
rect 20622 3720 20628 3732
rect 20220 3692 20628 3720
rect 20220 3680 20226 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 28960 3692 35894 3720
rect 28960 3680 28966 3692
rect 26206 3624 31708 3652
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 15703 3556 17969 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 17957 3553 17969 3556
rect 18003 3553 18015 3587
rect 19978 3584 19984 3596
rect 17957 3547 18015 3553
rect 18432 3556 19984 3584
rect 18432 3528 18460 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20806 3584 20812 3596
rect 20767 3556 20812 3584
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 22002 3544 22008 3596
rect 22060 3584 22066 3596
rect 26206 3584 26234 3624
rect 31570 3584 31576 3596
rect 22060 3556 26234 3584
rect 31531 3556 31576 3584
rect 22060 3544 22066 3556
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 31680 3584 31708 3624
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 35345 3655 35403 3661
rect 35345 3652 35357 3655
rect 31904 3624 35357 3652
rect 31904 3612 31910 3624
rect 35345 3621 35357 3624
rect 35391 3621 35403 3655
rect 35866 3652 35894 3692
rect 37366 3652 37372 3664
rect 35866 3624 37372 3652
rect 35345 3615 35403 3621
rect 37366 3612 37372 3624
rect 37424 3612 37430 3664
rect 36814 3584 36820 3596
rect 31680 3556 35894 3584
rect 36775 3556 36820 3584
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 14476 3488 16129 3516
rect 14369 3479 14427 3485
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 18414 3516 18420 3528
rect 18327 3488 18420 3516
rect 16117 3479 16175 3485
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20254 3516 20260 3528
rect 20211 3488 20260 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20625 3519 20683 3525
rect 20625 3485 20637 3519
rect 20671 3485 20683 3519
rect 31018 3516 31024 3528
rect 30979 3488 31024 3516
rect 20625 3479 20683 3485
rect 17770 3448 17776 3460
rect 17731 3420 17776 3448
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 20640 3448 20668 3479
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 33318 3516 33324 3528
rect 33279 3488 33324 3516
rect 33318 3476 33324 3488
rect 33376 3476 33382 3528
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 21726 3448 21732 3460
rect 20640 3420 21732 3448
rect 21726 3408 21732 3420
rect 21784 3408 21790 3460
rect 30834 3408 30840 3460
rect 30892 3448 30898 3460
rect 31205 3451 31263 3457
rect 31205 3448 31217 3451
rect 30892 3420 31217 3448
rect 30892 3408 30898 3420
rect 31205 3417 31217 3420
rect 31251 3417 31263 3451
rect 31205 3411 31263 3417
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 33980 3448 34008 3479
rect 31352 3420 34008 3448
rect 31352 3408 31358 3420
rect 34146 3408 34152 3460
rect 34204 3448 34210 3460
rect 35161 3451 35219 3457
rect 35161 3448 35173 3451
rect 34204 3420 35173 3448
rect 34204 3408 34210 3420
rect 35161 3417 35173 3420
rect 35207 3417 35219 3451
rect 35161 3411 35219 3417
rect 3568 3352 8984 3380
rect 18509 3383 18567 3389
rect 3568 3340 3574 3352
rect 18509 3349 18521 3383
rect 18555 3380 18567 3383
rect 19150 3380 19156 3392
rect 18555 3352 19156 3380
rect 18555 3349 18567 3352
rect 18509 3343 18567 3349
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19334 3380 19340 3392
rect 19295 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 23842 3380 23848 3392
rect 21968 3352 23848 3380
rect 21968 3340 21974 3352
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 32766 3340 32772 3392
rect 32824 3380 32830 3392
rect 33413 3383 33471 3389
rect 33413 3380 33425 3383
rect 32824 3352 33425 3380
rect 32824 3340 32830 3352
rect 33413 3349 33425 3352
rect 33459 3349 33471 3383
rect 33413 3343 33471 3349
rect 34057 3383 34115 3389
rect 34057 3349 34069 3383
rect 34103 3380 34115 3383
rect 34606 3380 34612 3392
rect 34103 3352 34612 3380
rect 34103 3349 34115 3352
rect 34057 3343 34115 3349
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 35866 3380 35894 3556
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 37826 3584 37832 3596
rect 37787 3556 37832 3584
rect 37826 3544 37832 3556
rect 37884 3544 37890 3596
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 37458 3408 37464 3460
rect 37516 3448 37522 3460
rect 38028 3448 38056 3479
rect 37516 3420 38056 3448
rect 37516 3408 37522 3420
rect 38654 3380 38660 3392
rect 35866 3352 38660 3380
rect 38654 3340 38660 3352
rect 38712 3340 38718 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2682 3176 2688 3188
rect 2643 3148 2688 3176
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 14366 3176 14372 3188
rect 3436 3148 14372 3176
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 2314 3040 2320 3052
rect 2179 3012 2320 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2406 3000 2412 3052
rect 2464 3040 2470 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2464 3012 2605 3040
rect 2464 3000 2470 3012
rect 2593 3009 2605 3012
rect 2639 3040 2651 3043
rect 3436 3040 3464 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 19242 3176 19248 3188
rect 17184 3148 19248 3176
rect 17184 3136 17190 3148
rect 19242 3136 19248 3148
rect 19300 3176 19306 3188
rect 30834 3176 30840 3188
rect 19300 3148 26234 3176
rect 30795 3148 30840 3176
rect 19300 3136 19306 3148
rect 3970 3068 3976 3120
rect 4028 3108 4034 3120
rect 7926 3108 7932 3120
rect 4028 3080 7932 3108
rect 4028 3068 4034 3080
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 19150 3108 19156 3120
rect 19111 3080 19156 3108
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 20714 3068 20720 3120
rect 20772 3108 20778 3120
rect 22005 3111 22063 3117
rect 22005 3108 22017 3111
rect 20772 3080 22017 3108
rect 20772 3068 20778 3080
rect 22005 3077 22017 3080
rect 22051 3077 22063 3111
rect 23658 3108 23664 3120
rect 23619 3080 23664 3108
rect 22005 3071 22063 3077
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 2639 3012 3464 3040
rect 5629 3043 5687 3049
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 3326 2972 3332 2984
rect 3287 2944 3332 2972
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 4982 2972 4988 2984
rect 4943 2944 4988 2972
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5644 2848 5672 3003
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 8662 3040 8668 3052
rect 5776 3012 5821 3040
rect 8623 3012 8668 3040
rect 5776 3000 5782 3012
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18969 3043 19027 3049
rect 18969 3040 18981 3043
rect 18564 3012 18981 3040
rect 18564 3000 18570 3012
rect 18969 3009 18981 3012
rect 19015 3009 19027 3043
rect 21818 3040 21824 3052
rect 21779 3012 21824 3040
rect 18969 3003 19027 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 26206 3040 26234 3148
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 35618 3176 35624 3188
rect 34900 3148 35624 3176
rect 32766 3108 32772 3120
rect 32727 3080 32772 3108
rect 32766 3068 32772 3080
rect 32824 3068 32830 3120
rect 30745 3043 30803 3049
rect 30745 3040 30757 3043
rect 26206 3012 30757 3040
rect 30745 3009 30757 3012
rect 30791 3040 30803 3043
rect 31294 3040 31300 3052
rect 30791 3012 31300 3040
rect 30791 3009 30803 3012
rect 30745 3003 30803 3009
rect 31294 3000 31300 3012
rect 31352 3000 31358 3052
rect 31389 3043 31447 3049
rect 31389 3009 31401 3043
rect 31435 3009 31447 3043
rect 32582 3040 32588 3052
rect 32543 3012 32588 3040
rect 31389 3003 31447 3009
rect 6362 2972 6368 2984
rect 6323 2944 6368 2972
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 6825 2935 6883 2941
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6840 2904 6868 2935
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 11514 2972 11520 2984
rect 11475 2944 11520 2972
rect 9125 2935 9183 2941
rect 5868 2876 6868 2904
rect 5868 2864 5874 2876
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9140 2904 9168 2935
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 14458 2972 14464 2984
rect 14419 2944 14464 2972
rect 11977 2935 12035 2941
rect 8444 2876 9168 2904
rect 8444 2864 8450 2876
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11992 2904 12020 2935
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14826 2972 14832 2984
rect 14787 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 16666 2972 16672 2984
rect 16627 2944 16672 2972
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16850 2972 16856 2984
rect 16811 2944 16856 2972
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 11020 2876 12020 2904
rect 11020 2864 11026 2876
rect 16758 2864 16764 2916
rect 16816 2904 16822 2916
rect 17144 2904 17172 2935
rect 18046 2932 18052 2984
rect 18104 2972 18110 2984
rect 19429 2975 19487 2981
rect 19429 2972 19441 2975
rect 18104 2944 19441 2972
rect 18104 2932 18110 2944
rect 19429 2941 19441 2944
rect 19475 2941 19487 2975
rect 31404 2972 31432 3003
rect 32582 3000 32588 3012
rect 32640 3000 32646 3052
rect 34900 3049 34928 3148
rect 35618 3136 35624 3148
rect 35676 3136 35682 3188
rect 35710 3136 35716 3188
rect 35768 3176 35774 3188
rect 37737 3179 37795 3185
rect 37737 3176 37749 3179
rect 35768 3148 37749 3176
rect 35768 3136 35774 3148
rect 37737 3145 37749 3148
rect 37783 3145 37795 3179
rect 37737 3139 37795 3145
rect 35069 3111 35127 3117
rect 35069 3077 35081 3111
rect 35115 3108 35127 3111
rect 35342 3108 35348 3120
rect 35115 3080 35348 3108
rect 35115 3077 35127 3080
rect 35069 3071 35127 3077
rect 35342 3068 35348 3080
rect 35400 3068 35406 3120
rect 38010 3108 38016 3120
rect 37971 3080 38016 3108
rect 38010 3068 38016 3080
rect 38068 3068 38074 3120
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 33318 2972 33324 2984
rect 31404 2944 33324 2972
rect 19429 2935 19487 2941
rect 33318 2932 33324 2944
rect 33376 2932 33382 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 35434 2972 35440 2984
rect 35395 2944 35440 2972
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 16816 2876 17172 2904
rect 16816 2864 16822 2876
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 1636 2808 2053 2836
rect 1636 2796 1642 2808
rect 2041 2805 2053 2808
rect 2087 2805 2099 2839
rect 5626 2836 5632 2848
rect 5539 2808 5632 2836
rect 2041 2799 2099 2805
rect 5626 2796 5632 2808
rect 5684 2836 5690 2848
rect 18322 2836 18328 2848
rect 5684 2808 18328 2836
rect 5684 2796 5690 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 31481 2839 31539 2845
rect 31481 2805 31493 2839
rect 31527 2836 31539 2839
rect 32490 2836 32496 2848
rect 31527 2808 32496 2836
rect 31527 2805 31539 2808
rect 31481 2799 31539 2805
rect 32490 2796 32496 2808
rect 32548 2796 32554 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5166 2632 5172 2644
rect 4755 2604 5172 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8846 2632 8852 2644
rect 8067 2604 8852 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 11698 2632 11704 2644
rect 10551 2604 11704 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 16117 2635 16175 2641
rect 16117 2601 16129 2635
rect 16163 2632 16175 2635
rect 16666 2632 16672 2644
rect 16163 2604 16672 2632
rect 16163 2601 16175 2604
rect 16117 2595 16175 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 16761 2635 16819 2641
rect 16761 2601 16773 2635
rect 16807 2632 16819 2635
rect 16850 2632 16856 2644
rect 16807 2604 16856 2632
rect 16807 2601 16819 2604
rect 16761 2595 16819 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17770 2632 17776 2644
rect 17451 2604 17776 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18601 2635 18659 2641
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 20070 2632 20076 2644
rect 18647 2604 20076 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21784 2604 21833 2632
rect 21784 2592 21790 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 31018 2632 31024 2644
rect 30979 2604 31024 2632
rect 21821 2595 21879 2601
rect 31018 2592 31024 2604
rect 31076 2592 31082 2644
rect 37458 2632 37464 2644
rect 37419 2604 37464 2632
rect 37458 2592 37464 2604
rect 37516 2592 37522 2644
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2564 4031 2567
rect 4982 2564 4988 2576
rect 4019 2536 4988 2564
rect 4019 2533 4031 2536
rect 3973 2527 4031 2533
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 5537 2567 5595 2573
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 6546 2564 6552 2576
rect 5583 2536 6552 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2564 10011 2567
rect 11514 2564 11520 2576
rect 9999 2536 11520 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 19334 2524 19340 2576
rect 19392 2524 19398 2576
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 19352 2496 19380 2524
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 19352 2468 19533 2496
rect 19521 2465 19533 2468
rect 19567 2465 19579 2499
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19521 2459 19579 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 32306 2496 32312 2508
rect 32267 2468 32312 2496
rect 32306 2456 32312 2468
rect 32364 2456 32370 2508
rect 32490 2496 32496 2508
rect 32451 2468 32496 2496
rect 32490 2456 32496 2468
rect 32548 2456 32554 2508
rect 32858 2496 32864 2508
rect 32819 2468 32864 2496
rect 32858 2456 32864 2468
rect 32916 2456 32922 2508
rect 34698 2496 34704 2508
rect 34659 2468 34704 2496
rect 34698 2456 34704 2468
rect 34756 2456 34762 2508
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4798 2428 4804 2440
rect 4111 2400 4804 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 7926 2428 7932 2440
rect 7887 2400 7932 2428
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 10410 2428 10416 2440
rect 10323 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16546 2400 16681 2428
rect 10428 2360 10456 2388
rect 16546 2360 16574 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 18414 2428 18420 2440
rect 17543 2400 18420 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 10428 2332 16574 2360
rect 16684 2292 16712 2391
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 19334 2428 19340 2440
rect 19295 2400 19340 2428
rect 19334 2388 19340 2400
rect 19392 2388 19398 2440
rect 18509 2363 18567 2369
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 18690 2360 18696 2372
rect 18555 2332 18696 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 34606 2320 34612 2372
rect 34664 2360 34670 2372
rect 34885 2363 34943 2369
rect 34885 2360 34897 2363
rect 34664 2332 34897 2360
rect 34664 2320 34670 2332
rect 34885 2329 34897 2332
rect 34931 2329 34943 2363
rect 34885 2323 34943 2329
rect 36541 2363 36599 2369
rect 36541 2329 36553 2363
rect 36587 2360 36599 2363
rect 37182 2360 37188 2372
rect 36587 2332 37188 2360
rect 36587 2329 36599 2332
rect 36541 2323 36599 2329
rect 37182 2320 37188 2332
rect 37240 2320 37246 2372
rect 20162 2292 20168 2304
rect 16684 2264 20168 2292
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 30006 1300 30012 1352
rect 30064 1340 30070 1352
rect 34514 1340 34520 1352
rect 30064 1312 34520 1340
rect 30064 1300 30070 1312
rect 34514 1300 34520 1312
rect 34572 1300 34578 1352
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 3424 37408 3476 37460
rect 7472 37408 7524 37460
rect 22468 37408 22520 37460
rect 36176 37408 36228 37460
rect 21824 37340 21876 37392
rect 23388 37340 23440 37392
rect 35348 37340 35400 37392
rect 11428 37272 11480 37324
rect 11704 37272 11756 37324
rect 15200 37315 15252 37324
rect 15200 37281 15209 37315
rect 15209 37281 15243 37315
rect 15243 37281 15252 37315
rect 15200 37272 15252 37281
rect 19984 37315 20036 37324
rect 19984 37281 19993 37315
rect 19993 37281 20027 37315
rect 20027 37281 20036 37315
rect 19984 37272 20036 37281
rect 22560 37272 22612 37324
rect 34796 37272 34848 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 2320 37247 2372 37256
rect 2320 37213 2329 37247
rect 2329 37213 2363 37247
rect 2363 37213 2372 37247
rect 2320 37204 2372 37213
rect 3424 37204 3476 37256
rect 6460 37204 6512 37256
rect 7748 37204 7800 37256
rect 9680 37204 9732 37256
rect 11520 37247 11572 37256
rect 11520 37213 11529 37247
rect 11529 37213 11563 37247
rect 11563 37213 11572 37247
rect 11520 37204 11572 37213
rect 14096 37247 14148 37256
rect 14096 37213 14105 37247
rect 14105 37213 14139 37247
rect 14139 37213 14148 37247
rect 14096 37204 14148 37213
rect 14832 37204 14884 37256
rect 17500 37204 17552 37256
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 20812 37204 20864 37256
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 7932 37136 7984 37188
rect 6736 37111 6788 37120
rect 6736 37077 6745 37111
rect 6745 37077 6779 37111
rect 6779 37077 6788 37111
rect 6736 37068 6788 37077
rect 10876 37136 10928 37188
rect 19984 37136 20036 37188
rect 22100 37136 22152 37188
rect 25872 37204 25924 37256
rect 28080 37247 28132 37256
rect 28080 37213 28089 37247
rect 28089 37213 28123 37247
rect 28123 37213 28132 37247
rect 28080 37204 28132 37213
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 33784 37204 33836 37256
rect 36728 37247 36780 37256
rect 36728 37213 36737 37247
rect 36737 37213 36771 37247
rect 36771 37213 36780 37247
rect 36728 37204 36780 37213
rect 36820 37204 36872 37256
rect 35348 37136 35400 37188
rect 12348 37068 12400 37120
rect 12440 37068 12492 37120
rect 17408 37068 17460 37120
rect 24308 37068 24360 37120
rect 24400 37111 24452 37120
rect 24400 37077 24409 37111
rect 24409 37077 24443 37111
rect 24443 37077 24452 37111
rect 24400 37068 24452 37077
rect 27896 37068 27948 37120
rect 37464 37111 37516 37120
rect 37464 37077 37473 37111
rect 37473 37077 37507 37111
rect 37507 37077 37516 37111
rect 37464 37068 37516 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 10876 36907 10928 36916
rect 10876 36873 10885 36907
rect 10885 36873 10919 36907
rect 10919 36873 10928 36907
rect 10876 36864 10928 36873
rect 12348 36864 12400 36916
rect 6736 36796 6788 36848
rect 20 36728 72 36780
rect 3424 36771 3476 36780
rect 3424 36737 3433 36771
rect 3433 36737 3467 36771
rect 3467 36737 3476 36771
rect 3424 36728 3476 36737
rect 3884 36660 3936 36712
rect 4160 36703 4212 36712
rect 4160 36669 4169 36703
rect 4169 36669 4203 36703
rect 4203 36669 4212 36703
rect 4160 36660 4212 36669
rect 7748 36592 7800 36644
rect 1860 36524 1912 36576
rect 3056 36524 3108 36576
rect 11520 36796 11572 36848
rect 10784 36771 10836 36780
rect 10784 36737 10793 36771
rect 10793 36737 10827 36771
rect 10827 36737 10836 36771
rect 10784 36728 10836 36737
rect 14096 36728 14148 36780
rect 17500 36771 17552 36780
rect 17500 36737 17509 36771
rect 17509 36737 17543 36771
rect 17543 36737 17552 36771
rect 17500 36728 17552 36737
rect 12256 36703 12308 36712
rect 12256 36669 12265 36703
rect 12265 36669 12299 36703
rect 12299 36669 12308 36703
rect 12256 36660 12308 36669
rect 12624 36660 12676 36712
rect 17684 36703 17736 36712
rect 17684 36669 17693 36703
rect 17693 36669 17727 36703
rect 17727 36669 17736 36703
rect 17684 36660 17736 36669
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 7932 36592 7984 36644
rect 12440 36592 12492 36644
rect 19984 36864 20036 36916
rect 21732 36864 21784 36916
rect 24400 36864 24452 36916
rect 24308 36839 24360 36848
rect 24308 36805 24317 36839
rect 24317 36805 24351 36839
rect 24351 36805 24360 36839
rect 24308 36796 24360 36805
rect 27896 36839 27948 36848
rect 27896 36805 27905 36839
rect 27905 36805 27939 36839
rect 27939 36805 27948 36839
rect 27896 36796 27948 36805
rect 37464 36796 37516 36848
rect 20812 36728 20864 36780
rect 21364 36728 21416 36780
rect 21824 36771 21876 36780
rect 21824 36737 21833 36771
rect 21833 36737 21867 36771
rect 21867 36737 21876 36771
rect 21824 36728 21876 36737
rect 23572 36728 23624 36780
rect 33784 36771 33836 36780
rect 33784 36737 33793 36771
rect 33793 36737 33827 36771
rect 33827 36737 33836 36771
rect 33784 36728 33836 36737
rect 34796 36728 34848 36780
rect 37188 36728 37240 36780
rect 20720 36660 20772 36712
rect 23020 36592 23072 36644
rect 23204 36592 23256 36644
rect 28540 36660 28592 36712
rect 29092 36703 29144 36712
rect 29092 36669 29101 36703
rect 29101 36669 29135 36703
rect 29135 36669 29144 36703
rect 29092 36660 29144 36669
rect 24676 36592 24728 36644
rect 21088 36524 21140 36576
rect 22376 36524 22428 36576
rect 36268 36524 36320 36576
rect 36452 36524 36504 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3884 36363 3936 36372
rect 3884 36329 3893 36363
rect 3893 36329 3927 36363
rect 3927 36329 3936 36363
rect 3884 36320 3936 36329
rect 7748 36320 7800 36372
rect 10784 36320 10836 36372
rect 12624 36363 12676 36372
rect 12624 36329 12633 36363
rect 12633 36329 12667 36363
rect 12667 36329 12676 36363
rect 12624 36320 12676 36329
rect 17684 36363 17736 36372
rect 17684 36329 17693 36363
rect 17693 36329 17727 36363
rect 17727 36329 17736 36363
rect 17684 36320 17736 36329
rect 19432 36320 19484 36372
rect 21364 36320 21416 36372
rect 24676 36320 24728 36372
rect 35348 36320 35400 36372
rect 2320 36252 2372 36304
rect 1308 36184 1360 36236
rect 3056 36227 3108 36236
rect 3056 36193 3065 36227
rect 3065 36193 3099 36227
rect 3099 36193 3108 36227
rect 3056 36184 3108 36193
rect 21272 36252 21324 36304
rect 7472 36184 7524 36236
rect 11428 36184 11480 36236
rect 22376 36227 22428 36236
rect 22376 36193 22385 36227
rect 22385 36193 22419 36227
rect 22419 36193 22428 36227
rect 22376 36184 22428 36193
rect 22560 36227 22612 36236
rect 22560 36193 22569 36227
rect 22569 36193 22603 36227
rect 22603 36193 22612 36227
rect 22560 36184 22612 36193
rect 36820 36252 36872 36304
rect 25872 36227 25924 36236
rect 25872 36193 25881 36227
rect 25881 36193 25915 36227
rect 25915 36193 25924 36227
rect 25872 36184 25924 36193
rect 26424 36227 26476 36236
rect 26424 36193 26433 36227
rect 26433 36193 26467 36227
rect 26467 36193 26476 36227
rect 26424 36184 26476 36193
rect 36268 36227 36320 36236
rect 36268 36193 36277 36227
rect 36277 36193 36311 36227
rect 36311 36193 36320 36227
rect 36268 36184 36320 36193
rect 36452 36227 36504 36236
rect 36452 36193 36461 36227
rect 36461 36193 36495 36227
rect 36495 36193 36504 36227
rect 36452 36184 36504 36193
rect 38108 36227 38160 36236
rect 38108 36193 38117 36227
rect 38117 36193 38151 36227
rect 38151 36193 38160 36227
rect 38108 36184 38160 36193
rect 12716 36159 12768 36168
rect 12716 36125 12725 36159
rect 12725 36125 12759 36159
rect 12759 36125 12768 36159
rect 12716 36116 12768 36125
rect 17316 36116 17368 36168
rect 23940 36116 23992 36168
rect 25228 36159 25280 36168
rect 25228 36125 25237 36159
rect 25237 36125 25271 36159
rect 25271 36125 25280 36159
rect 25228 36116 25280 36125
rect 34888 36116 34940 36168
rect 35440 36116 35492 36168
rect 35624 36159 35676 36168
rect 35624 36125 35633 36159
rect 35633 36125 35667 36159
rect 35667 36125 35676 36159
rect 35624 36116 35676 36125
rect 11888 36091 11940 36100
rect 11888 36057 11897 36091
rect 11897 36057 11931 36091
rect 11931 36057 11940 36091
rect 11888 36048 11940 36057
rect 21364 35980 21416 36032
rect 36452 35980 36504 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 11888 35776 11940 35828
rect 28356 35776 28408 35828
rect 29092 35776 29144 35828
rect 36728 35751 36780 35760
rect 36728 35717 36737 35751
rect 36737 35717 36771 35751
rect 36771 35717 36780 35751
rect 36728 35708 36780 35717
rect 12716 35640 12768 35692
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 34888 35683 34940 35692
rect 34888 35649 34897 35683
rect 34897 35649 34931 35683
rect 34931 35649 34940 35683
rect 34888 35640 34940 35649
rect 38016 35683 38068 35692
rect 38016 35649 38025 35683
rect 38025 35649 38059 35683
rect 38059 35649 38068 35683
rect 38016 35640 38068 35649
rect 24492 35572 24544 35624
rect 24584 35615 24636 35624
rect 24584 35581 24593 35615
rect 24593 35581 24627 35615
rect 24627 35581 24636 35615
rect 24584 35572 24636 35581
rect 35532 35572 35584 35624
rect 23296 35436 23348 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 24492 35275 24544 35284
rect 24492 35241 24501 35275
rect 24501 35241 24535 35275
rect 24535 35241 24544 35275
rect 24492 35232 24544 35241
rect 35532 35232 35584 35284
rect 36176 35096 36228 35148
rect 36452 35139 36504 35148
rect 36452 35105 36461 35139
rect 36461 35105 36495 35139
rect 36495 35105 36504 35139
rect 36452 35096 36504 35105
rect 38108 35139 38160 35148
rect 38108 35105 38117 35139
rect 38117 35105 38151 35139
rect 38151 35105 38160 35139
rect 38108 35096 38160 35105
rect 1584 35028 1636 35080
rect 24676 35028 24728 35080
rect 35440 35028 35492 35080
rect 37464 34892 37516 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 29276 34620 29328 34672
rect 32220 34620 32272 34672
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 27344 34552 27396 34604
rect 29644 34552 29696 34604
rect 37464 34595 37516 34604
rect 37464 34561 37473 34595
rect 37473 34561 37507 34595
rect 37507 34561 37516 34595
rect 37464 34552 37516 34561
rect 1768 34527 1820 34536
rect 1768 34493 1777 34527
rect 1777 34493 1811 34527
rect 1811 34493 1820 34527
rect 1768 34484 1820 34493
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 4620 34484 4672 34536
rect 5540 34484 5592 34536
rect 28264 34484 28316 34536
rect 30932 34484 30984 34536
rect 36452 34484 36504 34536
rect 36268 34348 36320 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1768 34144 1820 34196
rect 36268 34051 36320 34060
rect 36268 34017 36277 34051
rect 36277 34017 36311 34051
rect 36311 34017 36320 34051
rect 36268 34008 36320 34017
rect 36452 34051 36504 34060
rect 36452 34017 36461 34051
rect 36461 34017 36495 34051
rect 36495 34017 36504 34051
rect 36452 34008 36504 34017
rect 38108 34051 38160 34060
rect 38108 34017 38117 34051
rect 38117 34017 38151 34051
rect 38151 34017 38160 34051
rect 38108 34008 38160 34017
rect 17316 33940 17368 33992
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 29276 33532 29328 33584
rect 38016 33507 38068 33516
rect 38016 33473 38025 33507
rect 38025 33473 38059 33507
rect 38059 33473 38068 33507
rect 38016 33464 38068 33473
rect 24584 33439 24636 33448
rect 24584 33405 24593 33439
rect 24593 33405 24627 33439
rect 24627 33405 24636 33439
rect 24584 33396 24636 33405
rect 24768 33439 24820 33448
rect 24768 33405 24777 33439
rect 24777 33405 24811 33439
rect 24811 33405 24820 33439
rect 24768 33396 24820 33405
rect 37832 33371 37884 33380
rect 37832 33337 37841 33371
rect 37841 33337 37875 33371
rect 37875 33337 37884 33371
rect 37832 33328 37884 33337
rect 18604 33303 18656 33312
rect 18604 33269 18613 33303
rect 18613 33269 18647 33303
rect 18647 33269 18656 33303
rect 18604 33260 18656 33269
rect 36544 33303 36596 33312
rect 36544 33269 36553 33303
rect 36553 33269 36587 33303
rect 36587 33269 36596 33303
rect 36544 33260 36596 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 24584 33056 24636 33108
rect 3424 32784 3476 32836
rect 18604 32920 18656 32972
rect 36544 32920 36596 32972
rect 19156 32784 19208 32836
rect 36636 32784 36688 32836
rect 38108 32827 38160 32836
rect 38108 32793 38117 32827
rect 38117 32793 38151 32827
rect 38151 32793 38160 32827
rect 38108 32784 38160 32793
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 19156 32555 19208 32564
rect 19156 32521 19165 32555
rect 19165 32521 19199 32555
rect 19199 32521 19208 32555
rect 19156 32512 19208 32521
rect 24768 32512 24820 32564
rect 36636 32555 36688 32564
rect 36636 32521 36645 32555
rect 36645 32521 36679 32555
rect 36679 32521 36688 32555
rect 36636 32512 36688 32521
rect 20260 32376 20312 32428
rect 21272 32376 21324 32428
rect 12716 32308 12768 32360
rect 17224 32308 17276 32360
rect 37648 32376 37700 32428
rect 37924 32308 37976 32360
rect 1400 32172 1452 32224
rect 36268 32172 36320 32224
rect 36452 32172 36504 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 36268 31875 36320 31884
rect 36268 31841 36277 31875
rect 36277 31841 36311 31875
rect 36311 31841 36320 31875
rect 36268 31832 36320 31841
rect 36452 31875 36504 31884
rect 36452 31841 36461 31875
rect 36461 31841 36495 31875
rect 36495 31841 36504 31875
rect 36452 31832 36504 31841
rect 38108 31875 38160 31884
rect 38108 31841 38117 31875
rect 38117 31841 38151 31875
rect 38151 31841 38160 31875
rect 38108 31832 38160 31841
rect 36176 31764 36228 31816
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 2136 31331 2188 31340
rect 2136 31297 2145 31331
rect 2145 31297 2179 31331
rect 2179 31297 2188 31331
rect 2136 31288 2188 31297
rect 37464 31288 37516 31340
rect 35808 31263 35860 31272
rect 35808 31229 35817 31263
rect 35817 31229 35851 31263
rect 35851 31229 35860 31263
rect 35808 31220 35860 31229
rect 36176 31220 36228 31272
rect 9680 31084 9732 31136
rect 10968 31084 11020 31136
rect 38108 31127 38160 31136
rect 38108 31093 38117 31127
rect 38117 31093 38151 31127
rect 38151 31093 38160 31127
rect 38108 31084 38160 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 37372 30787 37424 30796
rect 37372 30753 37381 30787
rect 37381 30753 37415 30787
rect 37415 30753 37424 30787
rect 37372 30744 37424 30753
rect 4160 30719 4212 30728
rect 4160 30685 4169 30719
rect 4169 30685 4203 30719
rect 4203 30685 4212 30719
rect 4160 30676 4212 30685
rect 34888 30676 34940 30728
rect 37372 30608 37424 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4160 30268 4212 30320
rect 36728 30311 36780 30320
rect 34888 30243 34940 30252
rect 34888 30209 34897 30243
rect 34897 30209 34931 30243
rect 34931 30209 34940 30243
rect 34888 30200 34940 30209
rect 4620 30132 4672 30184
rect 5540 30175 5592 30184
rect 5540 30141 5549 30175
rect 5549 30141 5583 30175
rect 5583 30141 5592 30175
rect 5540 30132 5592 30141
rect 36728 30277 36737 30311
rect 36737 30277 36771 30311
rect 36771 30277 36780 30311
rect 36728 30268 36780 30277
rect 37372 30311 37424 30320
rect 37372 30277 37381 30311
rect 37381 30277 37415 30311
rect 37415 30277 37424 30311
rect 37372 30268 37424 30277
rect 37280 30243 37332 30252
rect 37280 30209 37289 30243
rect 37289 30209 37323 30243
rect 37323 30209 37332 30243
rect 37280 30200 37332 30209
rect 37924 30243 37976 30252
rect 37924 30209 37933 30243
rect 37933 30209 37967 30243
rect 37967 30209 37976 30243
rect 37924 30200 37976 30209
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4620 29792 4672 29844
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 37188 29699 37240 29708
rect 37188 29665 37197 29699
rect 37197 29665 37231 29699
rect 37231 29665 37240 29699
rect 37188 29656 37240 29665
rect 38108 29699 38160 29708
rect 38108 29665 38117 29699
rect 38117 29665 38151 29699
rect 38151 29665 38160 29699
rect 38108 29656 38160 29665
rect 4804 29588 4856 29640
rect 21732 29563 21784 29572
rect 21732 29529 21741 29563
rect 21741 29529 21775 29563
rect 21775 29529 21784 29563
rect 21732 29520 21784 29529
rect 37464 29520 37516 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 37464 29291 37516 29300
rect 37464 29257 37473 29291
rect 37473 29257 37507 29291
rect 37507 29257 37516 29291
rect 37464 29248 37516 29257
rect 37280 29112 37332 29164
rect 37464 29112 37516 29164
rect 37556 29044 37608 29096
rect 36452 28908 36504 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 21732 28704 21784 28756
rect 36452 28611 36504 28620
rect 36452 28577 36461 28611
rect 36461 28577 36495 28611
rect 36495 28577 36504 28611
rect 36452 28568 36504 28577
rect 38108 28611 38160 28620
rect 38108 28577 38117 28611
rect 38117 28577 38151 28611
rect 38151 28577 38160 28611
rect 38108 28568 38160 28577
rect 1768 28500 1820 28552
rect 8484 28500 8536 28552
rect 9772 28500 9824 28552
rect 18604 28500 18656 28552
rect 21824 28500 21876 28552
rect 32312 28543 32364 28552
rect 32312 28509 32321 28543
rect 32321 28509 32355 28543
rect 32355 28509 32364 28543
rect 32312 28500 32364 28509
rect 36268 28543 36320 28552
rect 36268 28509 36277 28543
rect 36277 28509 36311 28543
rect 36311 28509 36320 28543
rect 36268 28500 36320 28509
rect 21548 28475 21600 28484
rect 21548 28441 21557 28475
rect 21557 28441 21591 28475
rect 21591 28441 21600 28475
rect 21548 28432 21600 28441
rect 21916 28407 21968 28416
rect 21916 28373 21925 28407
rect 21925 28373 21959 28407
rect 21959 28373 21968 28407
rect 21916 28364 21968 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 19432 28092 19484 28144
rect 33324 28160 33376 28212
rect 1768 28067 1820 28076
rect 1768 28033 1777 28067
rect 1777 28033 1811 28067
rect 1811 28033 1820 28067
rect 1768 28024 1820 28033
rect 8484 28067 8536 28076
rect 8484 28033 8493 28067
rect 8493 28033 8527 28067
rect 8527 28033 8536 28067
rect 8484 28024 8536 28033
rect 18788 28067 18840 28076
rect 18788 28033 18797 28067
rect 18797 28033 18831 28067
rect 18831 28033 18840 28067
rect 18788 28024 18840 28033
rect 19340 28024 19392 28076
rect 1952 27999 2004 28008
rect 1952 27965 1961 27999
rect 1961 27965 1995 27999
rect 1995 27965 2004 27999
rect 1952 27956 2004 27965
rect 8668 27999 8720 28008
rect 1492 27888 1544 27940
rect 8668 27965 8677 27999
rect 8677 27965 8711 27999
rect 8711 27965 8720 27999
rect 8668 27956 8720 27965
rect 8300 27888 8352 27940
rect 18420 27956 18472 28008
rect 22468 28024 22520 28076
rect 31760 28024 31812 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 36268 28024 36320 28076
rect 22652 27999 22704 28008
rect 22652 27965 22661 27999
rect 22661 27965 22695 27999
rect 22695 27965 22704 27999
rect 32496 27999 32548 28008
rect 22652 27956 22704 27965
rect 32496 27965 32505 27999
rect 32505 27965 32539 27999
rect 32539 27965 32548 27999
rect 32496 27956 32548 27965
rect 32864 27999 32916 28008
rect 32864 27965 32873 27999
rect 32873 27965 32907 27999
rect 32907 27965 32916 27999
rect 32864 27956 32916 27965
rect 23296 27888 23348 27940
rect 23204 27820 23256 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1952 27616 2004 27668
rect 8668 27616 8720 27668
rect 32496 27616 32548 27668
rect 18604 27591 18656 27600
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 9772 27523 9824 27532
rect 9772 27489 9781 27523
rect 9781 27489 9815 27523
rect 9815 27489 9824 27523
rect 9772 27480 9824 27489
rect 9956 27480 10008 27532
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 18788 27548 18840 27600
rect 19432 27480 19484 27532
rect 20076 27548 20128 27600
rect 20628 27548 20680 27600
rect 28080 27548 28132 27600
rect 21824 27480 21876 27532
rect 22008 27523 22060 27532
rect 22008 27489 22017 27523
rect 22017 27489 22051 27523
rect 22051 27489 22060 27523
rect 22008 27480 22060 27489
rect 23296 27523 23348 27532
rect 23296 27489 23305 27523
rect 23305 27489 23339 27523
rect 23339 27489 23348 27523
rect 23296 27480 23348 27489
rect 9128 27455 9180 27464
rect 2228 27412 2280 27421
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 17408 27412 17460 27464
rect 17868 27412 17920 27464
rect 18328 27455 18380 27464
rect 18328 27421 18337 27455
rect 18337 27421 18371 27455
rect 18371 27421 18380 27455
rect 18328 27412 18380 27421
rect 18788 27412 18840 27464
rect 9956 27387 10008 27396
rect 9956 27353 9965 27387
rect 9965 27353 9999 27387
rect 9999 27353 10008 27387
rect 9956 27344 10008 27353
rect 10232 27276 10284 27328
rect 19340 27276 19392 27328
rect 20352 27276 20404 27328
rect 22652 27412 22704 27464
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 31760 27412 31812 27464
rect 22468 27344 22520 27396
rect 21732 27276 21784 27328
rect 22284 27276 22336 27328
rect 22928 27276 22980 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9956 27115 10008 27124
rect 9956 27081 9965 27115
rect 9965 27081 9999 27115
rect 9999 27081 10008 27115
rect 9956 27072 10008 27081
rect 10232 27072 10284 27124
rect 19432 27072 19484 27124
rect 21548 27072 21600 27124
rect 23020 27072 23072 27124
rect 18696 27004 18748 27056
rect 20076 27047 20128 27056
rect 20076 27013 20085 27047
rect 20085 27013 20119 27047
rect 20119 27013 20128 27047
rect 20076 27004 20128 27013
rect 20812 27004 20864 27056
rect 15200 26936 15252 26988
rect 18328 26936 18380 26988
rect 19340 26979 19392 26988
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 20536 26936 20588 26988
rect 17224 26911 17276 26920
rect 17224 26877 17233 26911
rect 17233 26877 17267 26911
rect 17267 26877 17276 26911
rect 17224 26868 17276 26877
rect 22008 26800 22060 26852
rect 10784 26732 10836 26784
rect 20076 26732 20128 26784
rect 22376 26732 22428 26784
rect 22928 26936 22980 26988
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 23388 26911 23440 26920
rect 23388 26877 23397 26911
rect 23397 26877 23431 26911
rect 23431 26877 23440 26911
rect 23388 26868 23440 26877
rect 38016 26979 38068 26988
rect 38016 26945 38025 26979
rect 38025 26945 38059 26979
rect 38059 26945 38068 26979
rect 38016 26936 38068 26945
rect 37280 26868 37332 26920
rect 22560 26732 22612 26784
rect 23204 26732 23256 26784
rect 23848 26732 23900 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18236 26528 18288 26580
rect 28080 26528 28132 26580
rect 2044 26392 2096 26444
rect 18236 26435 18288 26444
rect 18236 26401 18245 26435
rect 18245 26401 18279 26435
rect 18279 26401 18288 26435
rect 18236 26392 18288 26401
rect 19432 26392 19484 26444
rect 19984 26392 20036 26444
rect 1584 26324 1636 26376
rect 17500 26367 17552 26376
rect 17500 26333 17509 26367
rect 17509 26333 17543 26367
rect 17543 26333 17552 26367
rect 17500 26324 17552 26333
rect 18328 26324 18380 26376
rect 20536 26367 20588 26376
rect 20536 26333 20545 26367
rect 20545 26333 20579 26367
rect 20579 26333 20588 26367
rect 20536 26324 20588 26333
rect 21180 26324 21232 26376
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 22560 26367 22612 26376
rect 22560 26333 22569 26367
rect 22569 26333 22603 26367
rect 22603 26333 22612 26367
rect 22560 26324 22612 26333
rect 22744 26367 22796 26376
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 34704 26367 34756 26376
rect 34704 26333 34713 26367
rect 34713 26333 34747 26367
rect 34747 26333 34756 26367
rect 34704 26324 34756 26333
rect 36268 26367 36320 26376
rect 36268 26333 36277 26367
rect 36277 26333 36311 26367
rect 36311 26333 36320 26367
rect 36268 26324 36320 26333
rect 21088 26299 21140 26308
rect 21088 26265 21097 26299
rect 21097 26265 21131 26299
rect 21131 26265 21140 26299
rect 21088 26256 21140 26265
rect 21364 26256 21416 26308
rect 23296 26256 23348 26308
rect 37372 26256 37424 26308
rect 38200 26256 38252 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 22192 25984 22244 26036
rect 23020 25984 23072 26036
rect 23388 25984 23440 26036
rect 37372 26027 37424 26036
rect 3424 25959 3476 25968
rect 3424 25925 3433 25959
rect 3433 25925 3467 25959
rect 3467 25925 3476 25959
rect 3424 25916 3476 25925
rect 18420 25916 18472 25968
rect 37372 25993 37381 26027
rect 37381 25993 37415 26027
rect 37415 25993 37424 26027
rect 37372 25984 37424 25993
rect 23848 25959 23900 25968
rect 23848 25925 23857 25959
rect 23857 25925 23891 25959
rect 23891 25925 23900 25959
rect 23848 25916 23900 25925
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17500 25848 17552 25900
rect 20536 25891 20588 25900
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 21180 25848 21232 25900
rect 21916 25848 21968 25900
rect 22100 25848 22152 25900
rect 22376 25848 22428 25900
rect 33324 25848 33376 25900
rect 36268 25848 36320 25900
rect 37280 25891 37332 25900
rect 37280 25857 37289 25891
rect 37289 25857 37323 25891
rect 37323 25857 37332 25891
rect 37280 25848 37332 25857
rect 37924 25891 37976 25900
rect 37924 25857 37933 25891
rect 37933 25857 37967 25891
rect 37967 25857 37976 25891
rect 37924 25848 37976 25857
rect 2044 25780 2096 25832
rect 3516 25780 3568 25832
rect 20444 25780 20496 25832
rect 22652 25823 22704 25832
rect 22652 25789 22661 25823
rect 22661 25789 22695 25823
rect 22695 25789 22704 25823
rect 22652 25780 22704 25789
rect 34704 25780 34756 25832
rect 35808 25823 35860 25832
rect 35808 25789 35817 25823
rect 35817 25789 35851 25823
rect 35851 25789 35860 25823
rect 35808 25780 35860 25789
rect 37464 25712 37516 25764
rect 23480 25644 23532 25696
rect 24032 25687 24084 25696
rect 24032 25653 24041 25687
rect 24041 25653 24075 25687
rect 24075 25653 24084 25687
rect 24032 25644 24084 25653
rect 37924 25644 37976 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2044 25483 2096 25492
rect 2044 25449 2053 25483
rect 2053 25449 2087 25483
rect 2087 25449 2096 25483
rect 2044 25440 2096 25449
rect 21088 25440 21140 25492
rect 21548 25440 21600 25492
rect 22468 25440 22520 25492
rect 2320 25236 2372 25288
rect 18604 25279 18656 25288
rect 18604 25245 18613 25279
rect 18613 25245 18647 25279
rect 18647 25245 18656 25279
rect 18604 25236 18656 25245
rect 22376 25372 22428 25424
rect 20076 25347 20128 25356
rect 20076 25313 20085 25347
rect 20085 25313 20119 25347
rect 20119 25313 20128 25347
rect 20076 25304 20128 25313
rect 21732 25304 21784 25356
rect 22192 25236 22244 25288
rect 17960 25168 18012 25220
rect 21548 25211 21600 25220
rect 21548 25177 21557 25211
rect 21557 25177 21591 25211
rect 21591 25177 21600 25211
rect 21548 25168 21600 25177
rect 22468 25304 22520 25356
rect 22652 25440 22704 25492
rect 37832 25372 37884 25424
rect 28264 25304 28316 25356
rect 37924 25347 37976 25356
rect 37924 25313 37933 25347
rect 37933 25313 37967 25347
rect 37967 25313 37976 25347
rect 37924 25304 37976 25313
rect 22100 25100 22152 25152
rect 22468 25100 22520 25152
rect 22560 25100 22612 25152
rect 23020 25100 23072 25152
rect 23848 25236 23900 25288
rect 24308 25236 24360 25288
rect 38108 25279 38160 25288
rect 38108 25245 38117 25279
rect 38117 25245 38151 25279
rect 38151 25245 38160 25279
rect 38108 25236 38160 25245
rect 25872 25211 25924 25220
rect 25872 25177 25881 25211
rect 25881 25177 25915 25211
rect 25915 25177 25924 25211
rect 25872 25168 25924 25177
rect 36176 25168 36228 25220
rect 23572 25100 23624 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 24308 24939 24360 24948
rect 18604 24760 18656 24812
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 21088 24760 21140 24812
rect 21916 24803 21968 24812
rect 21916 24769 21926 24803
rect 21926 24769 21960 24803
rect 21960 24769 21968 24803
rect 21916 24760 21968 24769
rect 22100 24760 22152 24812
rect 23020 24828 23072 24880
rect 22468 24760 22520 24812
rect 23388 24803 23440 24812
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 4804 24624 4856 24676
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 24308 24905 24317 24939
rect 24317 24905 24351 24939
rect 24351 24905 24360 24939
rect 24308 24896 24360 24905
rect 25872 24939 25924 24948
rect 25872 24905 25881 24939
rect 25881 24905 25915 24939
rect 25915 24905 25924 24939
rect 25872 24896 25924 24905
rect 23572 24828 23624 24880
rect 23848 24760 23900 24812
rect 21272 24624 21324 24676
rect 23388 24624 23440 24676
rect 19064 24556 19116 24608
rect 21456 24556 21508 24608
rect 21916 24556 21968 24608
rect 23204 24556 23256 24608
rect 23756 24624 23808 24676
rect 25596 24760 25648 24812
rect 38108 24760 38160 24812
rect 23664 24556 23716 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1860 24148 1912 24200
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 18604 24216 18656 24268
rect 21364 24352 21416 24404
rect 22560 24352 22612 24404
rect 21916 24284 21968 24336
rect 22836 24284 22888 24336
rect 20352 24191 20404 24200
rect 18788 24080 18840 24132
rect 20352 24157 20361 24191
rect 20361 24157 20395 24191
rect 20395 24157 20404 24191
rect 20352 24148 20404 24157
rect 20536 24148 20588 24200
rect 20904 24148 20956 24200
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 22100 24148 22152 24200
rect 22652 24148 22704 24200
rect 23204 24148 23256 24200
rect 23388 24259 23440 24268
rect 23388 24225 23398 24259
rect 23398 24225 23432 24259
rect 23432 24225 23440 24259
rect 23388 24216 23440 24225
rect 24400 24327 24452 24336
rect 24400 24293 24409 24327
rect 24409 24293 24443 24327
rect 24443 24293 24452 24327
rect 24400 24284 24452 24293
rect 25504 24259 25556 24268
rect 25504 24225 25513 24259
rect 25513 24225 25547 24259
rect 25547 24225 25556 24259
rect 25504 24216 25556 24225
rect 27344 24259 27396 24268
rect 27344 24225 27353 24259
rect 27353 24225 27387 24259
rect 27387 24225 27396 24259
rect 27344 24216 27396 24225
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 21364 24012 21416 24064
rect 21824 24012 21876 24064
rect 23112 24012 23164 24064
rect 23296 24080 23348 24132
rect 38108 24148 38160 24200
rect 23848 24080 23900 24132
rect 25688 24123 25740 24132
rect 25688 24089 25697 24123
rect 25697 24089 25731 24123
rect 25731 24089 25740 24123
rect 25688 24080 25740 24089
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 21088 23851 21140 23860
rect 21088 23817 21097 23851
rect 21097 23817 21131 23851
rect 21131 23817 21140 23851
rect 21088 23808 21140 23817
rect 21364 23808 21416 23860
rect 25688 23851 25740 23860
rect 3700 23783 3752 23792
rect 3700 23749 3709 23783
rect 3709 23749 3743 23783
rect 3743 23749 3752 23783
rect 3700 23740 3752 23749
rect 18420 23783 18472 23792
rect 18420 23749 18429 23783
rect 18429 23749 18463 23783
rect 18463 23749 18472 23783
rect 18420 23740 18472 23749
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 17224 23672 17276 23724
rect 17868 23672 17920 23724
rect 2044 23647 2096 23656
rect 2044 23613 2053 23647
rect 2053 23613 2087 23647
rect 2087 23613 2096 23647
rect 2044 23604 2096 23613
rect 18604 23672 18656 23724
rect 19432 23672 19484 23724
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 20536 23604 20588 23656
rect 22652 23672 22704 23724
rect 22836 23740 22888 23792
rect 28172 23740 28224 23792
rect 23112 23672 23164 23724
rect 24400 23672 24452 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 37280 23715 37332 23724
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 22744 23604 22796 23656
rect 18604 23536 18656 23588
rect 18788 23536 18840 23588
rect 20352 23536 20404 23588
rect 23296 23536 23348 23588
rect 21456 23468 21508 23520
rect 22928 23468 22980 23520
rect 25504 23468 25556 23520
rect 37924 23468 37976 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2044 23264 2096 23316
rect 23296 23264 23348 23316
rect 28080 23264 28132 23316
rect 35532 23264 35584 23316
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 6552 23060 6604 23112
rect 19432 23060 19484 23112
rect 17316 22992 17368 23044
rect 19340 22992 19392 23044
rect 35624 23196 35676 23248
rect 37280 23196 37332 23248
rect 37188 23171 37240 23180
rect 37188 23137 37197 23171
rect 37197 23137 37231 23171
rect 37231 23137 37240 23171
rect 37188 23128 37240 23137
rect 37924 23171 37976 23180
rect 37924 23137 37933 23171
rect 37933 23137 37967 23171
rect 37967 23137 37976 23171
rect 37924 23128 37976 23137
rect 38108 23171 38160 23180
rect 38108 23137 38117 23171
rect 38117 23137 38151 23171
rect 38151 23137 38160 23171
rect 38108 23128 38160 23137
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22100 23060 22152 23112
rect 24584 23060 24636 23112
rect 28080 23060 28132 23112
rect 21180 22992 21232 23044
rect 20996 22924 21048 22976
rect 22100 22924 22152 22976
rect 28356 22924 28408 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 20720 22763 20772 22772
rect 20720 22729 20729 22763
rect 20729 22729 20763 22763
rect 20763 22729 20772 22763
rect 20720 22720 20772 22729
rect 25596 22720 25648 22772
rect 20904 22652 20956 22704
rect 19432 22627 19484 22636
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 19708 22584 19760 22636
rect 21088 22584 21140 22636
rect 21916 22584 21968 22636
rect 23480 22652 23532 22704
rect 28356 22695 28408 22704
rect 28356 22661 28365 22695
rect 28365 22661 28399 22695
rect 28399 22661 28408 22695
rect 28356 22652 28408 22661
rect 22560 22584 22612 22636
rect 28172 22627 28224 22636
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 28172 22584 28224 22593
rect 37740 22584 37792 22636
rect 20260 22516 20312 22568
rect 30012 22559 30064 22568
rect 30012 22525 30021 22559
rect 30021 22525 30055 22559
rect 30055 22525 30064 22559
rect 30012 22516 30064 22525
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 22468 22380 22520 22432
rect 36544 22423 36596 22432
rect 36544 22389 36553 22423
rect 36553 22389 36587 22423
rect 36587 22389 36596 22423
rect 36544 22380 36596 22389
rect 36636 22380 36688 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 21824 22108 21876 22160
rect 23848 22176 23900 22228
rect 23480 22040 23532 22092
rect 24032 22040 24084 22092
rect 36544 22040 36596 22092
rect 38108 22083 38160 22092
rect 38108 22049 38117 22083
rect 38117 22049 38151 22083
rect 38151 22049 38160 22083
rect 38108 22040 38160 22049
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 22008 22015 22060 22024
rect 22008 21981 22050 22015
rect 22050 21981 22060 22015
rect 22008 21972 22060 21981
rect 19432 21947 19484 21956
rect 19432 21913 19441 21947
rect 19441 21913 19475 21947
rect 19475 21913 19484 21947
rect 19432 21904 19484 21913
rect 36636 21904 36688 21956
rect 22008 21836 22060 21888
rect 22192 21836 22244 21888
rect 23572 21836 23624 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 19432 21496 19484 21548
rect 20260 21496 20312 21548
rect 22192 21496 22244 21548
rect 23480 21496 23532 21548
rect 31760 21496 31812 21548
rect 37648 21496 37700 21548
rect 21916 21471 21968 21480
rect 21916 21437 21925 21471
rect 21925 21437 21959 21471
rect 21959 21437 21968 21471
rect 21916 21428 21968 21437
rect 23388 21403 23440 21412
rect 23388 21369 23397 21403
rect 23397 21369 23431 21403
rect 23431 21369 23440 21403
rect 23388 21360 23440 21369
rect 19800 21335 19852 21344
rect 19800 21301 19809 21335
rect 19809 21301 19843 21335
rect 19843 21301 19852 21335
rect 19800 21292 19852 21301
rect 19984 21292 20036 21344
rect 20444 21292 20496 21344
rect 36268 21292 36320 21344
rect 36636 21292 36688 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 20352 21020 20404 21072
rect 20168 20952 20220 21004
rect 22008 20952 22060 21004
rect 22468 20927 22520 20936
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 36268 20995 36320 21004
rect 36268 20961 36277 20995
rect 36277 20961 36311 20995
rect 36311 20961 36320 20995
rect 36268 20952 36320 20961
rect 36636 20952 36688 21004
rect 38108 20995 38160 21004
rect 38108 20961 38117 20995
rect 38117 20961 38151 20995
rect 38151 20961 38160 20995
rect 38108 20952 38160 20961
rect 31760 20884 31812 20936
rect 19800 20816 19852 20868
rect 34520 20816 34572 20868
rect 23204 20748 23256 20800
rect 24216 20748 24268 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 22928 20544 22980 20596
rect 23204 20587 23256 20596
rect 23204 20553 23213 20587
rect 23213 20553 23247 20587
rect 23247 20553 23256 20587
rect 23204 20544 23256 20553
rect 2136 20476 2188 20528
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 22100 20476 22152 20528
rect 23388 20519 23440 20528
rect 23388 20485 23397 20519
rect 23397 20485 23431 20519
rect 23431 20485 23440 20519
rect 23388 20476 23440 20485
rect 24216 20519 24268 20528
rect 24216 20485 24225 20519
rect 24225 20485 24259 20519
rect 24259 20485 24268 20519
rect 24216 20476 24268 20485
rect 21180 20408 21232 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 18604 20340 18656 20392
rect 25872 20383 25924 20392
rect 25872 20349 25881 20383
rect 25881 20349 25915 20383
rect 25915 20349 25924 20383
rect 25872 20340 25924 20349
rect 21364 20272 21416 20324
rect 1676 20204 1728 20256
rect 2136 20247 2188 20256
rect 2136 20213 2145 20247
rect 2145 20213 2179 20247
rect 2179 20213 2188 20247
rect 2136 20204 2188 20213
rect 2780 20247 2832 20256
rect 2780 20213 2789 20247
rect 2789 20213 2823 20247
rect 2823 20213 2832 20247
rect 2780 20204 2832 20213
rect 22192 20204 22244 20256
rect 37924 20204 37976 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2136 19932 2188 19984
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 22100 19932 22152 19984
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 23204 19864 23256 19916
rect 37188 19907 37240 19916
rect 37188 19873 37197 19907
rect 37197 19873 37231 19907
rect 37231 19873 37240 19907
rect 37188 19864 37240 19873
rect 37924 19907 37976 19916
rect 37924 19873 37933 19907
rect 37933 19873 37967 19907
rect 37967 19873 37976 19907
rect 37924 19864 37976 19873
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 31760 19839 31812 19848
rect 31760 19805 31769 19839
rect 31769 19805 31803 19839
rect 31803 19805 31812 19839
rect 31760 19796 31812 19805
rect 38108 19839 38160 19848
rect 38108 19805 38117 19839
rect 38117 19805 38151 19839
rect 38151 19805 38160 19839
rect 38108 19796 38160 19805
rect 23848 19771 23900 19780
rect 23848 19737 23857 19771
rect 23857 19737 23891 19771
rect 23891 19737 23900 19771
rect 23848 19728 23900 19737
rect 24584 19771 24636 19780
rect 24584 19737 24593 19771
rect 24593 19737 24627 19771
rect 24627 19737 24636 19771
rect 24584 19728 24636 19737
rect 35624 19728 35676 19780
rect 22100 19660 22152 19712
rect 32312 19660 32364 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 24584 19456 24636 19508
rect 2780 19388 2832 19440
rect 22008 19388 22060 19440
rect 32312 19431 32364 19440
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 23940 19363 23992 19372
rect 23940 19329 23949 19363
rect 23949 19329 23983 19363
rect 23983 19329 23992 19363
rect 23940 19320 23992 19329
rect 32312 19397 32321 19431
rect 32321 19397 32355 19431
rect 32355 19397 32364 19431
rect 32312 19388 32364 19397
rect 38108 19320 38160 19372
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 31760 19184 31812 19236
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1400 18912 1452 18964
rect 12440 18776 12492 18828
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 22284 18411 22336 18420
rect 22284 18377 22293 18411
rect 22293 18377 22327 18411
rect 22327 18377 22336 18411
rect 22284 18368 22336 18377
rect 20720 18232 20772 18284
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 27252 18028 27304 18080
rect 27620 18071 27672 18080
rect 27620 18037 27629 18071
rect 27629 18037 27663 18071
rect 27663 18037 27672 18071
rect 27620 18028 27672 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17688 1636 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 27620 17756 27672 17808
rect 2780 17688 2832 17697
rect 27252 17731 27304 17740
rect 27252 17697 27261 17731
rect 27261 17697 27295 17731
rect 27295 17697 27304 17731
rect 27252 17688 27304 17697
rect 1952 17552 2004 17604
rect 28908 17595 28960 17604
rect 28908 17561 28917 17595
rect 28917 17561 28951 17595
rect 28951 17561 28960 17595
rect 28908 17552 28960 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 9128 17144 9180 17196
rect 20628 17144 20680 17196
rect 29552 17076 29604 17128
rect 34520 17076 34572 17128
rect 3608 16983 3660 16992
rect 3608 16949 3617 16983
rect 3617 16949 3651 16983
rect 3651 16949 3660 16983
rect 3608 16940 3660 16949
rect 38108 16940 38160 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 29552 16779 29604 16788
rect 29552 16745 29561 16779
rect 29561 16745 29595 16779
rect 29595 16745 29604 16779
rect 29552 16736 29604 16745
rect 3424 16532 3476 16584
rect 20628 16668 20680 16720
rect 19340 16600 19392 16652
rect 37648 16643 37700 16652
rect 37648 16609 37657 16643
rect 37657 16609 37691 16643
rect 37691 16609 37700 16643
rect 37648 16600 37700 16609
rect 38108 16643 38160 16652
rect 38108 16609 38117 16643
rect 38117 16609 38151 16643
rect 38151 16609 38160 16643
rect 38108 16600 38160 16609
rect 37556 16464 37608 16516
rect 3240 16396 3292 16448
rect 4068 16396 4120 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 37556 16235 37608 16244
rect 37556 16201 37565 16235
rect 37565 16201 37599 16235
rect 37599 16201 37608 16235
rect 37556 16192 37608 16201
rect 3240 16167 3292 16176
rect 3240 16133 3249 16167
rect 3249 16133 3283 16167
rect 3283 16133 3292 16167
rect 3240 16124 3292 16133
rect 4068 16167 4120 16176
rect 4068 16133 4077 16167
rect 4077 16133 4111 16167
rect 4111 16133 4120 16167
rect 4068 16124 4120 16133
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 3608 16056 3660 16108
rect 19064 16056 19116 16108
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 3424 15920 3476 15972
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4436 15512 4488 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 19064 15512 19116 15564
rect 38108 15444 38160 15496
rect 21824 15376 21876 15428
rect 4252 15308 4304 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4252 15079 4304 15088
rect 4252 15045 4261 15079
rect 4261 15045 4295 15079
rect 4295 15045 4304 15079
rect 4252 15036 4304 15045
rect 2136 14968 2188 15020
rect 4436 15011 4488 15020
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 17960 14968 18012 15020
rect 37648 14968 37700 15020
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 3056 14764 3108 14816
rect 19800 14807 19852 14816
rect 19800 14773 19809 14807
rect 19809 14773 19843 14807
rect 19843 14773 19852 14807
rect 19800 14764 19852 14773
rect 37924 14764 37976 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 19800 14467 19852 14476
rect 19800 14433 19809 14467
rect 19809 14433 19843 14467
rect 19843 14433 19852 14467
rect 19800 14424 19852 14433
rect 37188 14467 37240 14476
rect 37188 14433 37197 14467
rect 37197 14433 37231 14467
rect 37231 14433 37240 14467
rect 37188 14424 37240 14433
rect 37924 14467 37976 14476
rect 37924 14433 37933 14467
rect 37933 14433 37967 14467
rect 37967 14433 37976 14467
rect 37924 14424 37976 14433
rect 38108 14467 38160 14476
rect 38108 14433 38117 14467
rect 38117 14433 38151 14467
rect 38151 14433 38160 14467
rect 38108 14424 38160 14433
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 19432 14288 19484 14340
rect 34520 14288 34572 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 18696 13880 18748 13932
rect 19432 13880 19484 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 37832 13719 37884 13728
rect 37832 13685 37841 13719
rect 37841 13685 37875 13719
rect 37875 13685 37884 13719
rect 37832 13676 37884 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3516 13472 3568 13524
rect 37188 13379 37240 13388
rect 37188 13345 37197 13379
rect 37197 13345 37231 13379
rect 37231 13345 37240 13379
rect 37188 13336 37240 13345
rect 37832 13336 37884 13388
rect 1400 13268 1452 13320
rect 37556 13200 37608 13252
rect 3976 13132 4028 13184
rect 19432 13132 19484 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 37556 12971 37608 12980
rect 37556 12937 37565 12971
rect 37565 12937 37599 12971
rect 37599 12937 37608 12971
rect 37556 12928 37608 12937
rect 2228 12792 2280 12844
rect 3700 12792 3752 12844
rect 20260 12792 20312 12844
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 37740 12792 37792 12844
rect 1584 12588 1636 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 37188 12291 37240 12300
rect 37188 12257 37197 12291
rect 37197 12257 37231 12291
rect 37231 12257 37240 12291
rect 37188 12248 37240 12257
rect 35808 12180 35860 12232
rect 37280 12112 37332 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 37832 11704 37884 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2044 11636 2096 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 36268 11500 36320 11552
rect 37648 11543 37700 11552
rect 37648 11509 37657 11543
rect 37657 11509 37691 11543
rect 37691 11509 37700 11543
rect 37648 11500 37700 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 35808 11339 35860 11348
rect 35808 11305 35817 11339
rect 35817 11305 35851 11339
rect 35851 11305 35860 11339
rect 35808 11296 35860 11305
rect 36268 11203 36320 11212
rect 36268 11169 36277 11203
rect 36277 11169 36311 11203
rect 36311 11169 36320 11203
rect 36268 11160 36320 11169
rect 37648 11160 37700 11212
rect 38108 11203 38160 11212
rect 38108 11169 38117 11203
rect 38117 11169 38151 11203
rect 38151 11169 38160 11203
rect 38108 11160 38160 11169
rect 2688 11092 2740 11144
rect 18144 11092 18196 11144
rect 18512 11092 18564 11144
rect 20168 11092 20220 11144
rect 20260 11067 20312 11076
rect 20260 11033 20269 11067
rect 20269 11033 20303 11067
rect 20303 11033 20312 11067
rect 20260 11024 20312 11033
rect 37832 11024 37884 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 37280 10752 37332 10804
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 20260 10616 20312 10668
rect 37832 10616 37884 10668
rect 6092 10412 6144 10464
rect 36268 10412 36320 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6276 10072 6328 10124
rect 36268 10115 36320 10124
rect 36268 10081 36277 10115
rect 36277 10081 36311 10115
rect 36311 10081 36320 10115
rect 36268 10072 36320 10081
rect 38108 10115 38160 10124
rect 38108 10081 38117 10115
rect 38117 10081 38151 10115
rect 38151 10081 38160 10115
rect 38108 10072 38160 10081
rect 36452 9979 36504 9988
rect 36452 9945 36461 9979
rect 36461 9945 36495 9979
rect 36495 9945 36504 9979
rect 36452 9936 36504 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 36452 9664 36504 9716
rect 18420 9528 18472 9580
rect 37372 9571 37424 9580
rect 37372 9537 37381 9571
rect 37381 9537 37415 9571
rect 37415 9537 37424 9571
rect 37372 9528 37424 9537
rect 1400 9324 1452 9376
rect 37924 9324 37976 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 37188 9027 37240 9036
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 37924 9027 37976 9036
rect 37924 8993 37933 9027
rect 37933 8993 37967 9027
rect 37967 8993 37976 9027
rect 37924 8984 37976 8993
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 1952 8848 2004 8900
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2136 8440 2188 8492
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 19340 8440 19392 8492
rect 38108 8440 38160 8492
rect 4160 8372 4212 8424
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 3056 8304 3108 8356
rect 8300 8304 8352 8356
rect 3240 8236 3292 8288
rect 20628 8236 20680 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8300 8032 8352 8084
rect 9588 8032 9640 8084
rect 3056 7939 3108 7948
rect 3056 7905 3065 7939
rect 3065 7905 3099 7939
rect 3099 7905 3108 7939
rect 3056 7896 3108 7905
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 22008 7939 22060 7948
rect 22008 7905 22017 7939
rect 22017 7905 22051 7939
rect 22051 7905 22060 7939
rect 22008 7896 22060 7905
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 18604 7828 18656 7880
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 1400 7803 1452 7812
rect 1400 7769 1409 7803
rect 1409 7769 1443 7803
rect 1443 7769 1452 7803
rect 1400 7760 1452 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 20444 7352 20496 7404
rect 9404 7148 9456 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 9772 6672 9824 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 1952 6196 2004 6248
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2136 5652 2188 5704
rect 2412 5652 2464 5704
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3332 5312 3384 5364
rect 23940 5312 23992 5364
rect 10416 4972 10468 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 38108 4972 38160 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9680 4700 9732 4752
rect 3240 4632 3292 4684
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 37188 4675 37240 4684
rect 2872 4564 2924 4616
rect 18512 4564 18564 4616
rect 37188 4641 37197 4675
rect 37197 4641 37231 4675
rect 37231 4641 37240 4675
rect 37188 4632 37240 4641
rect 38108 4675 38160 4684
rect 38108 4641 38117 4675
rect 38117 4641 38151 4675
rect 38151 4641 38160 4675
rect 38108 4632 38160 4641
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20260 4564 20312 4616
rect 10600 4539 10652 4548
rect 10600 4505 10609 4539
rect 10609 4505 10643 4539
rect 10643 4505 10652 4539
rect 10600 4496 10652 4505
rect 37924 4539 37976 4548
rect 37924 4505 37933 4539
rect 37933 4505 37967 4539
rect 37967 4505 37976 4539
rect 37924 4496 37976 4505
rect 17960 4428 18012 4480
rect 20812 4471 20864 4480
rect 20812 4437 20821 4471
rect 20821 4437 20855 4471
rect 20855 4437 20864 4471
rect 20812 4428 20864 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 10600 4224 10652 4276
rect 37924 4224 37976 4276
rect 3516 4156 3568 4208
rect 17960 4199 18012 4208
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 3884 4020 3936 4072
rect 17960 4165 17969 4199
rect 17969 4165 18003 4199
rect 18003 4165 18012 4199
rect 17960 4156 18012 4165
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 22560 4088 22612 4140
rect 31852 4088 31904 4140
rect 3332 3952 3384 4004
rect 23664 3952 23716 4004
rect 34520 4020 34572 4072
rect 37280 4088 37332 4140
rect 37740 4020 37792 4072
rect 1400 3884 1452 3936
rect 6460 3884 6512 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9312 3884 9364 3936
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 22284 3884 22336 3936
rect 35716 3952 35768 4004
rect 32312 3927 32364 3936
rect 32312 3893 32321 3927
rect 32321 3893 32355 3927
rect 32355 3893 32364 3927
rect 32312 3884 32364 3893
rect 32588 3884 32640 3936
rect 34704 3884 34756 3936
rect 35348 3884 35400 3936
rect 35624 3927 35676 3936
rect 35624 3893 35633 3927
rect 35633 3893 35667 3927
rect 35667 3893 35676 3927
rect 35624 3884 35676 3893
rect 37832 3884 37884 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 664 3612 716 3664
rect 2872 3544 2924 3596
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 8668 3476 8720 3528
rect 2688 3408 2740 3460
rect 4620 3451 4672 3460
rect 4620 3417 4629 3451
rect 4629 3417 4663 3451
rect 4663 3417 4672 3451
rect 4620 3408 4672 3417
rect 5724 3408 5776 3460
rect 3516 3340 3568 3392
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 14280 3476 14332 3528
rect 20168 3680 20220 3732
rect 20628 3680 20680 3732
rect 28908 3680 28960 3732
rect 19984 3544 20036 3596
rect 20812 3587 20864 3596
rect 20812 3553 20821 3587
rect 20821 3553 20855 3587
rect 20855 3553 20864 3587
rect 20812 3544 20864 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 22008 3544 22060 3596
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 31852 3612 31904 3664
rect 37372 3612 37424 3664
rect 36820 3587 36872 3596
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 20260 3476 20312 3528
rect 31024 3519 31076 3528
rect 17776 3451 17828 3460
rect 17776 3417 17785 3451
rect 17785 3417 17819 3451
rect 17819 3417 17828 3451
rect 17776 3408 17828 3417
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 33324 3519 33376 3528
rect 33324 3485 33333 3519
rect 33333 3485 33367 3519
rect 33367 3485 33376 3519
rect 33324 3476 33376 3485
rect 21732 3408 21784 3460
rect 30840 3408 30892 3460
rect 31300 3408 31352 3460
rect 34152 3408 34204 3460
rect 19156 3340 19208 3392
rect 19340 3383 19392 3392
rect 19340 3349 19349 3383
rect 19349 3349 19383 3383
rect 19383 3349 19392 3383
rect 19340 3340 19392 3349
rect 21916 3340 21968 3392
rect 23848 3340 23900 3392
rect 32772 3340 32824 3392
rect 34612 3340 34664 3392
rect 36820 3553 36829 3587
rect 36829 3553 36863 3587
rect 36863 3553 36872 3587
rect 36820 3544 36872 3553
rect 37832 3587 37884 3596
rect 37832 3553 37841 3587
rect 37841 3553 37875 3587
rect 37875 3553 37884 3587
rect 37832 3544 37884 3553
rect 37464 3408 37516 3460
rect 38660 3340 38712 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 2320 3000 2372 3052
rect 2412 3000 2464 3052
rect 14372 3136 14424 3188
rect 17132 3136 17184 3188
rect 19248 3136 19300 3188
rect 30840 3179 30892 3188
rect 3976 3068 4028 3120
rect 7932 3068 7984 3120
rect 19156 3111 19208 3120
rect 19156 3077 19165 3111
rect 19165 3077 19199 3111
rect 19199 3077 19208 3111
rect 19156 3068 19208 3077
rect 20720 3068 20772 3120
rect 23664 3111 23716 3120
rect 23664 3077 23673 3111
rect 23673 3077 23707 3111
rect 23707 3077 23716 3111
rect 23664 3068 23716 3077
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 8668 3043 8720 3052
rect 5724 3000 5776 3009
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 18512 3000 18564 3052
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 30840 3145 30849 3179
rect 30849 3145 30883 3179
rect 30883 3145 30892 3179
rect 30840 3136 30892 3145
rect 32772 3111 32824 3120
rect 32772 3077 32781 3111
rect 32781 3077 32815 3111
rect 32815 3077 32824 3111
rect 32772 3068 32824 3077
rect 31300 3000 31352 3052
rect 32588 3043 32640 3052
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 8852 2975 8904 2984
rect 5816 2864 5868 2916
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 11520 2975 11572 2984
rect 8392 2864 8444 2916
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 14464 2975 14516 2984
rect 10968 2864 11020 2916
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 16856 2975 16908 2984
rect 16856 2941 16865 2975
rect 16865 2941 16899 2975
rect 16899 2941 16908 2975
rect 16856 2932 16908 2941
rect 16764 2864 16816 2916
rect 18052 2932 18104 2984
rect 32588 3009 32597 3043
rect 32597 3009 32631 3043
rect 32631 3009 32640 3043
rect 32588 3000 32640 3009
rect 35624 3136 35676 3188
rect 35716 3136 35768 3188
rect 35348 3068 35400 3120
rect 38016 3111 38068 3120
rect 38016 3077 38025 3111
rect 38025 3077 38059 3111
rect 38059 3077 38068 3111
rect 38016 3068 38068 3077
rect 33324 2932 33376 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 35440 2975 35492 2984
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 1584 2796 1636 2848
rect 5632 2796 5684 2848
rect 18328 2796 18380 2848
rect 32496 2796 32548 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5172 2592 5224 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 8852 2592 8904 2644
rect 11704 2592 11756 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 16672 2592 16724 2644
rect 16856 2592 16908 2644
rect 17776 2592 17828 2644
rect 20076 2592 20128 2644
rect 21732 2592 21784 2644
rect 31024 2635 31076 2644
rect 31024 2601 31033 2635
rect 31033 2601 31067 2635
rect 31067 2601 31076 2635
rect 31024 2592 31076 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 4988 2524 5040 2576
rect 6552 2524 6604 2576
rect 11520 2524 11572 2576
rect 19340 2524 19392 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 32312 2499 32364 2508
rect 32312 2465 32321 2499
rect 32321 2465 32355 2499
rect 32355 2465 32364 2499
rect 32312 2456 32364 2465
rect 32496 2499 32548 2508
rect 32496 2465 32505 2499
rect 32505 2465 32539 2499
rect 32539 2465 32548 2499
rect 32496 2456 32548 2465
rect 32864 2499 32916 2508
rect 32864 2465 32873 2499
rect 32873 2465 32907 2499
rect 32907 2465 32916 2499
rect 32864 2456 32916 2465
rect 34704 2499 34756 2508
rect 34704 2465 34713 2499
rect 34713 2465 34747 2499
rect 34747 2465 34756 2499
rect 34704 2456 34756 2465
rect 4804 2388 4856 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 18420 2388 18472 2440
rect 19340 2431 19392 2440
rect 19340 2397 19349 2431
rect 19349 2397 19383 2431
rect 19383 2397 19392 2431
rect 19340 2388 19392 2397
rect 18696 2320 18748 2372
rect 34612 2320 34664 2372
rect 37188 2320 37240 2372
rect 20168 2252 20220 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 30012 1300 30064 1352
rect 34520 1300 34572 1352
<< metal2 >>
rect -10 39200 102 40000
rect 634 39200 746 40000
rect 1278 39200 1390 40000
rect 1922 39200 2034 40000
rect 2566 39200 2678 40000
rect 3854 39200 3966 40000
rect 4498 39200 4610 40000
rect 5142 39200 5254 40000
rect 5786 39200 5898 40000
rect 6430 39200 6542 40000
rect 7074 39200 7186 40000
rect 7718 39200 7830 40000
rect 8312 39222 8892 39250
rect 32 36786 60 39200
rect 20 36780 72 36786
rect 20 36722 72 36728
rect 1320 36242 1348 39200
rect 1964 37618 1992 39200
rect 3330 38856 3386 38865
rect 3330 38791 3386 38800
rect 1504 37590 1992 37618
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 36825 1440 37198
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1308 36236 1360 36242
rect 1308 36178 1360 36184
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1504 27946 1532 37590
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 1860 36576 1912 36582
rect 1860 36518 1912 36524
rect 1872 35894 1900 36518
rect 2332 36310 2360 37198
rect 3056 36576 3108 36582
rect 3056 36518 3108 36524
rect 2320 36304 2372 36310
rect 2320 36246 2372 36252
rect 3068 36242 3096 36518
rect 3056 36236 3108 36242
rect 3056 36178 3108 36184
rect 1872 35866 2084 35894
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1596 34610 1624 35022
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 1780 34202 1808 34478
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1780 28082 1808 28494
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1952 28008 2004 28014
rect 1952 27950 2004 27956
rect 1492 27940 1544 27946
rect 1492 27882 1544 27888
rect 1964 27674 1992 27950
rect 1952 27668 2004 27674
rect 1952 27610 2004 27616
rect 2056 26450 2084 35866
rect 2778 34776 2834 34785
rect 2778 34711 2834 34720
rect 2792 34542 2820 34711
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 25906 1624 26318
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 2044 25832 2096 25838
rect 2044 25774 2096 25780
rect 2056 25498 2084 25774
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1872 23730 1900 24142
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 2044 23656 2096 23662
rect 2044 23598 2096 23604
rect 2056 23322 2084 23598
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1872 23118 1900 23151
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 2148 20534 2176 31282
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2136 20528 2188 20534
rect 2136 20470 2188 20476
rect 2240 20466 2268 27406
rect 3344 26234 3372 38791
rect 3422 37496 3478 37505
rect 3422 37431 3424 37440
rect 3476 37431 3478 37440
rect 3424 37402 3476 37408
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3436 36786 3464 37198
rect 3896 36802 3924 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 3424 36780 3476 36786
rect 3896 36774 4200 36802
rect 3424 36722 3476 36728
rect 4172 36718 4200 36774
rect 3884 36712 3936 36718
rect 3884 36654 3936 36660
rect 4160 36712 4212 36718
rect 4160 36654 4212 36660
rect 3896 36378 3924 36654
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 3884 36372 3936 36378
rect 3884 36314 3936 36320
rect 3698 36136 3754 36145
rect 3698 36071 3754 36080
rect 3422 33416 3478 33425
rect 3422 33351 3478 33360
rect 3436 32842 3464 33351
rect 3424 32836 3476 32842
rect 3424 32778 3476 32784
rect 3344 26206 3464 26234
rect 3436 25974 3464 26206
rect 3424 25968 3476 25974
rect 3424 25910 3476 25916
rect 3514 25936 3570 25945
rect 3514 25871 3570 25880
rect 3528 25838 3556 25871
rect 3516 25832 3568 25838
rect 3516 25774 3568 25780
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 18970 1440 19790
rect 1688 19378 1716 20198
rect 2148 19990 2176 20198
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19825 1900 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2148 19145 2176 19246
rect 2134 19136 2190 19145
rect 2134 19071 2190 19080
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17746 1624 18022
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1964 17338 1992 17546
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16574 2084 17138
rect 2056 16546 2176 16574
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15745 1624 15982
rect 1582 15736 1638 15745
rect 1582 15671 1638 15680
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 2148 15026 2176 16546
rect 1398 14991 1454 15000
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1400 14408 1452 14414
rect 1398 14376 1400 14385
rect 1452 14376 1454 14385
rect 1398 14311 1454 14320
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13705 1900 13806
rect 1858 13696 1914 13705
rect 1858 13631 1914 13640
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12306 1440 13262
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12306 1624 12582
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1688 10674 1716 11630
rect 2056 11354 2084 11630
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9042 1440 9318
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 8945 1900 8978
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2148 8498 2176 14962
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 1412 7585 1440 7754
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 2240 6914 2268 12786
rect 2148 6886 2268 6914
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6322 1624 6734
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1952 6248 2004 6254
rect 2044 6248 2096 6254
rect 1952 6190 2004 6196
rect 2042 6216 2044 6225
rect 2096 6216 2098 6225
rect 1964 5914 1992 6190
rect 2042 6151 2098 6160
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2148 5710 2176 6886
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 676 800 704 3606
rect 1412 2514 1440 3878
rect 2332 3058 2360 25230
rect 3712 23798 3740 36071
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4632 34542 4660 37726
rect 6472 37262 6500 39200
rect 7472 37460 7524 37466
rect 7472 37402 7524 37408
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6748 36854 6776 37062
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 7484 36242 7512 37402
rect 7760 37262 7788 39200
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 7932 37188 7984 37194
rect 7932 37130 7984 37136
rect 7944 36650 7972 37130
rect 7748 36644 7800 36650
rect 7748 36586 7800 36592
rect 7932 36644 7984 36650
rect 7932 36586 7984 36592
rect 7760 36378 7788 36586
rect 7748 36372 7800 36378
rect 7748 36314 7800 36320
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 5540 34536 5592 34542
rect 5540 34478 5592 34484
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4160 30728 4212 30734
rect 4160 30670 4212 30676
rect 4172 30326 4200 30670
rect 4160 30320 4212 30326
rect 4160 30262 4212 30268
rect 5552 30190 5580 34478
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29850 4660 30126
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4816 24682 4844 29582
rect 8312 27946 8340 39222
rect 8864 39114 8892 39222
rect 9006 39200 9118 40000
rect 9650 39200 9762 40000
rect 9968 39222 10180 39250
rect 9048 39114 9076 39200
rect 8864 39086 9076 39114
rect 9692 37262 9720 39200
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 8484 28552 8536 28558
rect 8484 28494 8536 28500
rect 8496 28082 8524 28494
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8668 28008 8720 28014
rect 8668 27950 8720 27956
rect 8300 27940 8352 27946
rect 8300 27882 8352 27888
rect 8680 27674 8708 27950
rect 8668 27668 8720 27674
rect 8668 27610 8720 27616
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2792 19446 2820 20198
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 16182 3280 16390
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3436 16114 3464 16526
rect 3620 16114 3648 16934
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16182 4108 16390
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 8498 2728 11086
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2884 6914 2912 14894
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14482 3096 14758
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 7954 3096 8298
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 7954 3280 8230
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 2792 6886 2912 6914
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 3058 2452 5646
rect 2792 3618 2820 6886
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2884 4146 2912 4558
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2608 3590 2820 3618
rect 3252 3602 3280 4626
rect 3344 4185 3372 5306
rect 3330 4176 3386 4185
rect 3330 4111 3386 4120
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 2872 3596 2924 3602
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2514 1624 2790
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2608 800 2636 3590
rect 2872 3538 2924 3544
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2700 3194 2728 3402
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2792 2514 2820 2751
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2884 2145 2912 3538
rect 3344 3074 3372 3946
rect 3252 3046 3372 3074
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 3252 800 3280 3046
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3344 1465 3372 2926
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3436 762 3464 15914
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15094 4292 15302
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4448 15026 4476 15506
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3528 13530 3556 13806
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3712 12850 3740 13806
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3514 4856 3570 4865
rect 3514 4791 3570 4800
rect 3528 4214 3556 4791
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3738 3924 4014
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3534 4016 13126
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4160 8424 4212 8430
rect 4080 8372 4160 8378
rect 4080 8366 4212 8372
rect 4080 8350 4200 8366
rect 4080 8265 4108 8350
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3976 3528 4028 3534
rect 3514 3496 3570 3505
rect 3976 3470 4028 3476
rect 3514 3431 3570 3440
rect 3528 3398 3556 3431
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3988 3126 4016 3470
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 1714 4660 3402
rect 4816 2446 4844 24618
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6564 10674 6592 23054
rect 9140 17202 9168 27406
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10130 6132 10406
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5736 3058 5764 3402
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5000 2582 5028 2926
rect 5184 2650 5212 2926
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 5644 2446 5672 2790
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 4540 1686 4660 1714
rect 3712 870 3924 898
rect 3712 762 3740 870
rect 3896 800 3924 870
rect 4540 800 4568 1686
rect 5828 800 5856 2858
rect 6288 1170 6316 10066
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 8090 8340 8298
rect 9600 8090 9628 8366
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7410 9168 7822
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 6866 9444 7142
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9692 4758 9720 31078
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9784 27538 9812 28494
rect 9968 27538 9996 39222
rect 10152 39114 10180 39222
rect 10294 39200 10406 40000
rect 10938 39200 11050 40000
rect 11582 39200 11694 40000
rect 12226 39200 12338 40000
rect 12870 39200 12982 40000
rect 14158 39200 14270 40000
rect 14802 39200 14914 40000
rect 15446 39200 15558 40000
rect 16090 39200 16202 40000
rect 16734 39200 16846 40000
rect 17378 39200 17490 40000
rect 18022 39200 18134 40000
rect 19310 39200 19422 40000
rect 19954 39200 20066 40000
rect 20598 39200 20710 40000
rect 21242 39200 21354 40000
rect 21886 39200 21998 40000
rect 22530 39200 22642 40000
rect 23174 39200 23286 40000
rect 24462 39200 24574 40000
rect 25106 39200 25218 40000
rect 25750 39200 25862 40000
rect 26394 39200 26506 40000
rect 27038 39200 27150 40000
rect 27682 39200 27794 40000
rect 28326 39200 28438 40000
rect 29614 39200 29726 40000
rect 30258 39200 30370 40000
rect 30902 39200 31014 40000
rect 31546 39200 31658 40000
rect 32190 39200 32302 40000
rect 32834 39200 32946 40000
rect 33478 39200 33590 40000
rect 34766 39200 34878 40000
rect 35410 39200 35522 40000
rect 36054 39200 36166 40000
rect 36698 39200 36810 40000
rect 37342 39200 37454 40000
rect 37986 39200 38098 40000
rect 38630 39200 38742 40000
rect 39274 39200 39386 40000
rect 10336 39114 10364 39200
rect 10152 39086 10364 39114
rect 10876 37188 10928 37194
rect 10876 37130 10928 37136
rect 10888 36922 10916 37130
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 10784 36780 10836 36786
rect 10784 36722 10836 36728
rect 10796 36378 10824 36722
rect 10784 36372 10836 36378
rect 10784 36314 10836 36320
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9956 27396 10008 27402
rect 9956 27338 10008 27344
rect 9968 27130 9996 27338
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10244 27130 10272 27270
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10796 26790 10824 36314
rect 10980 31142 11008 39200
rect 11624 37346 11652 39200
rect 11624 37330 11744 37346
rect 11428 37324 11480 37330
rect 11624 37324 11756 37330
rect 11624 37318 11704 37324
rect 11428 37266 11480 37272
rect 11704 37266 11756 37272
rect 11440 36242 11468 37266
rect 11520 37256 11572 37262
rect 11520 37198 11572 37204
rect 11532 36854 11560 37198
rect 11520 36848 11572 36854
rect 11520 36790 11572 36796
rect 12268 36718 12296 39200
rect 14844 37262 14872 39200
rect 15200 37324 15252 37330
rect 15200 37266 15252 37272
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 12440 37120 12492 37126
rect 12440 37062 12492 37068
rect 12360 36922 12388 37062
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12256 36712 12308 36718
rect 12256 36654 12308 36660
rect 12452 36650 12480 37062
rect 14108 36786 14136 37198
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12440 36644 12492 36650
rect 12440 36586 12492 36592
rect 12636 36378 12664 36654
rect 12624 36372 12676 36378
rect 12624 36314 12676 36320
rect 11428 36236 11480 36242
rect 11428 36178 11480 36184
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 11888 36100 11940 36106
rect 11888 36042 11940 36048
rect 11900 35834 11928 36042
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 12728 35698 12756 36110
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12728 32366 12756 35634
rect 12716 32360 12768 32366
rect 12716 32302 12768 32308
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 15212 26994 15240 37266
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17328 33998 17356 36110
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 17236 26926 17264 32302
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 16574 12480 18770
rect 12452 16546 13584 16574
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6730 9812 7142
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 6472 3602 6500 3878
rect 9140 3602 9168 3878
rect 9324 3602 9352 3878
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6380 2650 6408 2926
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6564 2582 6592 2926
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 7944 2446 7972 3062
rect 8680 3058 8708 3470
rect 9876 3346 9904 6802
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4690 10456 4966
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10612 4282 10640 4490
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9692 3318 9904 3346
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 6288 1142 6500 1170
rect 6472 800 6500 1142
rect 8404 800 8432 2858
rect 8864 2650 8892 2926
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9692 800 9720 3318
rect 10428 2446 10456 4082
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10980 800 11008 2858
rect 11532 2582 11560 2926
rect 11716 2650 11744 2926
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 13556 800 13584 16546
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3058 14320 3470
rect 17144 3194 17172 25842
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17236 23730 17264 24142
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17328 23050 17356 33934
rect 17420 27470 17448 37062
rect 17512 36786 17540 37198
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 18064 36718 18092 39200
rect 19996 37330 20024 39200
rect 19984 37324 20036 37330
rect 19984 37266 20036 37272
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 17684 36712 17736 36718
rect 17684 36654 17736 36660
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 17696 36378 17724 36654
rect 19444 36378 19472 37198
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36922 20024 37130
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 20640 36802 20668 39200
rect 20812 37256 20864 37262
rect 20812 37198 20864 37204
rect 20640 36774 20760 36802
rect 20824 36786 20852 37198
rect 20732 36718 20760 36774
rect 20812 36780 20864 36786
rect 20812 36722 20864 36728
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 17684 36372 17736 36378
rect 17684 36314 17736 36320
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18616 32978 18644 33254
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 32570 19196 32778
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19156 32564 19208 32570
rect 19156 32506 19208 32512
rect 20260 32428 20312 32434
rect 20260 32370 20312 32376
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17512 25906 17540 26318
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17880 23730 17908 27406
rect 18340 26994 18368 27406
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 18248 26450 18276 26522
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18248 26234 18276 26386
rect 18340 26382 18368 26930
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18156 26206 18276 26234
rect 17960 25220 18012 25226
rect 17960 25162 18012 25168
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17972 15026 18000 25162
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18156 11150 18184 26206
rect 18432 25974 18460 27950
rect 18616 27606 18644 28494
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 18800 27606 18828 28018
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18788 27600 18840 27606
rect 18788 27542 18840 27548
rect 18616 26234 18644 27542
rect 18800 27470 18828 27542
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 19352 27334 19380 28018
rect 19444 27538 19472 28086
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18524 26206 18644 26234
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18418 24168 18474 24177
rect 18418 24103 18474 24112
rect 18432 23798 18460 24103
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18432 9586 18460 23734
rect 18524 11150 18552 26206
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18616 24818 18644 25230
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18616 24274 18644 24754
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18616 23730 18644 24210
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18616 20398 18644 23530
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 6914 18460 9522
rect 18616 7886 18644 20334
rect 18708 13938 18736 26998
rect 19352 26994 19380 27270
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19444 26450 19472 27066
rect 20088 27062 20116 27542
rect 20076 27056 20128 27062
rect 20076 26998 20128 27004
rect 20088 26790 20116 26998
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19076 24614 19104 24686
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 18786 24304 18842 24313
rect 18786 24239 18842 24248
rect 18800 24138 18828 24239
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18800 23594 18828 24074
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 19076 16114 19104 24550
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23118 19472 23666
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19352 16658 19380 22986
rect 19444 22642 19472 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19720 22030 19748 22578
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19444 21554 19472 21898
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19996 21434 20024 26386
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 19444 21406 20024 21434
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19076 15570 19104 16050
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19444 14498 19472 21406
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19812 20874 19840 21286
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19352 14470 19472 14498
rect 19812 14482 19840 14758
rect 19800 14476 19852 14482
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 19352 8498 19380 14470
rect 19800 14418 19852 14424
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19444 14074 19472 14282
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13190 19472 13874
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 18340 6886 18460 6914
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4146 17816 4966
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 4214 18000 4422
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14384 2446 14412 3130
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 14476 2650 14504 2926
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14844 800 14872 2926
rect 16684 2650 16712 2926
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16776 800 16804 2858
rect 16868 2650 16896 2926
rect 17788 2650 17816 3402
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18064 800 18092 2926
rect 18340 2854 18368 6886
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18432 2446 18460 3470
rect 18524 3058 18552 4558
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19168 3126 19196 3334
rect 19260 3194 19288 3470
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 19352 2582 19380 3334
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 19340 2440 19392 2446
rect 19444 2394 19472 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 3602 20024 21286
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20088 2650 20116 25298
rect 20272 22574 20300 32370
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20364 24206 20392 27270
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20548 26382 20576 26930
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20548 25906 20576 26318
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20364 23594 20392 24142
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 21010 20208 21966
rect 20272 21706 20300 22510
rect 20272 21678 20392 21706
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20272 12850 20300 21490
rect 20364 21078 20392 21678
rect 20456 21350 20484 25774
rect 20534 24848 20590 24857
rect 20534 24783 20536 24792
rect 20588 24783 20590 24792
rect 20536 24754 20588 24760
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20548 23662 20576 24142
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20352 21072 20404 21078
rect 20352 21014 20404 21020
rect 20640 17202 20668 27542
rect 20824 27062 20852 36722
rect 21088 36576 21140 36582
rect 21088 36518 21140 36524
rect 21100 35894 21128 36518
rect 21284 36310 21312 39200
rect 21824 37392 21876 37398
rect 21824 37334 21876 37340
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 21376 36378 21404 36722
rect 21364 36372 21416 36378
rect 21364 36314 21416 36320
rect 21272 36304 21324 36310
rect 21272 36246 21324 36252
rect 21376 36038 21404 36314
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21376 35894 21404 35974
rect 21744 35894 21772 36858
rect 21836 36786 21864 37334
rect 21928 37210 21956 39200
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 21928 37194 22140 37210
rect 21928 37188 22152 37194
rect 21928 37182 22100 37188
rect 22100 37130 22152 37136
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22388 36242 22416 36518
rect 22376 36236 22428 36242
rect 22376 36178 22428 36184
rect 21100 35866 21220 35894
rect 21376 35866 21496 35894
rect 21744 35866 21864 35894
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 21192 26382 21220 35866
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 21100 25498 21128 26250
rect 21192 25906 21220 26318
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21284 24834 21312 32370
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21192 24806 21312 24834
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20732 18766 20760 22714
rect 20916 22710 20944 24142
rect 21100 23866 21128 24754
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 21008 22982 21036 23666
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 21100 22642 21128 23802
rect 21192 23050 21220 24806
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24206 21312 24618
rect 21376 24410 21404 26250
rect 21468 24614 21496 35866
rect 21732 29572 21784 29578
rect 21732 29514 21784 29520
rect 21744 28762 21772 29514
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21836 28558 21864 35866
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21548 28484 21600 28490
rect 21548 28426 21600 28432
rect 21560 27130 21588 28426
rect 21836 27538 21864 28494
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 21732 27328 21784 27334
rect 21732 27270 21784 27276
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 25226 21588 25434
rect 21744 25362 21772 27270
rect 21928 26024 21956 28358
rect 22480 28082 22508 37402
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 22572 36242 22600 37266
rect 23216 36650 23244 39200
rect 23388 37392 23440 37398
rect 23388 37334 23440 37340
rect 23020 36644 23072 36650
rect 23020 36586 23072 36592
rect 23204 36644 23256 36650
rect 23204 36586 23256 36592
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22020 26858 22048 27474
rect 22480 27402 22508 28018
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22664 27470 22692 27950
rect 23032 27470 23060 36586
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23308 27946 23336 35430
rect 23400 29714 23428 37334
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23584 36786 23612 37198
rect 24308 37120 24360 37126
rect 24308 37062 24360 37068
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24320 36854 24348 37062
rect 24412 36922 24440 37062
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24308 36848 24360 36854
rect 24308 36790 24360 36796
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23940 36168 23992 36174
rect 23940 36110 23992 36116
rect 23952 35698 23980 36110
rect 24504 35894 24532 39200
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 24676 36644 24728 36650
rect 24676 36586 24728 36592
rect 24688 36378 24716 36586
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 25884 36242 25912 37198
rect 26436 36242 26464 39200
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 27896 37120 27948 37126
rect 27896 37062 27948 37068
rect 27908 36854 27936 37062
rect 27896 36848 27948 36854
rect 27896 36790 27948 36796
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 26424 36236 26476 36242
rect 26424 36178 26476 36184
rect 25228 36168 25280 36174
rect 25228 36110 25280 36116
rect 24504 35866 24624 35894
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 24596 35630 24624 35866
rect 24492 35624 24544 35630
rect 24492 35566 24544 35572
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24504 35290 24532 35566
rect 24492 35284 24544 35290
rect 24492 35226 24544 35232
rect 24676 35080 24728 35086
rect 24676 35022 24728 35028
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24596 33114 24624 33390
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23296 27940 23348 27946
rect 23296 27882 23348 27888
rect 23204 27872 23256 27878
rect 23204 27814 23256 27820
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 22296 26382 22324 27270
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22192 26036 22244 26042
rect 21928 25996 22048 26024
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21732 25356 21784 25362
rect 21732 25298 21784 25304
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21928 24818 21956 25842
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21928 24342 21956 24550
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21272 24200 21324 24206
rect 22020 24188 22048 25996
rect 22192 25978 22244 25984
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25158 22140 25842
rect 22204 25294 22232 25978
rect 22388 25906 22416 26726
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22388 25430 22416 25842
rect 22480 25498 22508 27338
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22940 26994 22968 27270
rect 23032 27130 23060 27406
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 26382 22600 26726
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22664 25498 22692 25774
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 22376 25424 22428 25430
rect 22376 25366 22428 25372
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22112 24818 22140 25094
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22100 24200 22152 24206
rect 22020 24160 22100 24188
rect 21272 24142 21324 24148
rect 22100 24142 22152 24148
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21376 23866 21404 24006
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21192 20466 21220 22986
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21376 19854 21404 20266
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21468 19666 21496 23462
rect 21836 23118 21864 24006
rect 22112 23730 22140 24142
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 23118 22140 23666
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21928 22522 21956 22578
rect 21836 22494 21956 22522
rect 21836 22166 21864 22494
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21376 19638 21496 19666
rect 21376 18766 21404 19638
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 20732 18290 20760 18702
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20640 16726 20668 17138
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 21836 15434 21864 22102
rect 22020 22030 22048 22374
rect 22008 22024 22060 22030
rect 21928 21972 22008 21978
rect 21928 21966 22060 21972
rect 21928 21950 22048 21966
rect 21928 21486 21956 21950
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 22020 21010 22048 21830
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22112 20534 22140 22918
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21554 22232 21830
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22020 19446 22048 20402
rect 22112 19990 22140 20470
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22204 19922 22232 20198
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 22112 19378 22140 19654
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 18426 22324 19246
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20180 6914 20208 11086
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20272 10674 20300 11018
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7954 20668 8230
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7410 20484 7822
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20180 6886 20300 6914
rect 20272 4622 20300 6886
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19392 2388 19472 2394
rect 19340 2382 19472 2388
rect 18696 2372 18748 2378
rect 19352 2366 19472 2382
rect 18696 2314 18748 2320
rect 18708 800 18736 2314
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2450
rect 20180 2310 20208 3674
rect 20272 3534 20300 4558
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3738 20668 4082
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20732 3126 20760 3878
rect 20824 3602 20852 4422
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 21284 800 21312 3538
rect 21732 3460 21784 3466
rect 21732 3402 21784 3408
rect 21744 2650 21772 3402
rect 21836 3058 21864 3878
rect 22020 3602 22048 7890
rect 22388 6914 22416 25366
rect 22480 25362 22508 25434
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22480 24818 22508 25094
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22572 24698 22600 25094
rect 22480 24670 22600 24698
rect 22480 22522 22508 24670
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22572 22642 22600 24346
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22664 23730 22692 24142
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22756 23662 22784 26318
rect 23032 26042 23060 27066
rect 23216 26994 23244 27814
rect 23308 27538 23336 27882
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23020 26036 23072 26042
rect 23020 25978 23072 25984
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 24886 23060 25094
rect 23020 24880 23072 24886
rect 23020 24822 23072 24828
rect 23216 24614 23244 26726
rect 23400 26382 23428 26862
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 26308 23348 26314
rect 23296 26250 23348 26256
rect 23204 24608 23256 24614
rect 23124 24568 23204 24596
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22848 23798 22876 24278
rect 23124 24070 23152 24568
rect 23204 24550 23256 24556
rect 23308 24290 23336 26250
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23400 24818 23428 25978
rect 23860 25974 23888 26726
rect 23848 25968 23900 25974
rect 23848 25910 23900 25916
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23492 25242 23520 25638
rect 23860 25294 23888 25910
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 23848 25288 23900 25294
rect 23492 25214 23796 25242
rect 23848 25230 23900 25236
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 23216 24262 23336 24290
rect 23400 24274 23428 24618
rect 23388 24268 23440 24274
rect 23216 24206 23244 24262
rect 23388 24210 23440 24216
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 22836 23792 22888 23798
rect 22836 23734 22888 23740
rect 23124 23730 23152 24006
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 23308 23594 23336 24074
rect 23296 23588 23348 23594
rect 23296 23530 23348 23536
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22480 22494 22600 22522
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 20942 22508 22374
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22572 19334 22600 22494
rect 22940 20602 22968 23462
rect 23308 23322 23336 23530
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23492 22710 23520 25214
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24886 23612 25094
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23492 21554 23520 22034
rect 23584 21894 23612 24822
rect 23768 24682 23796 25214
rect 23860 24818 23888 25230
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23756 24676 23808 24682
rect 23756 24618 23808 24624
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23676 24206 23704 24550
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23860 22234 23888 24074
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 24044 22098 24072 25638
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 24320 24954 24348 25230
rect 24308 24948 24360 24954
rect 24308 24890 24360 24896
rect 24400 24336 24452 24342
rect 24688 24313 24716 35022
rect 24768 33448 24820 33454
rect 24768 33390 24820 33396
rect 24780 32570 24808 33390
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24400 24278 24452 24284
rect 24674 24304 24730 24313
rect 24412 23730 24440 24278
rect 24674 24239 24730 24248
rect 25240 24177 25268 36110
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 25872 25220 25924 25226
rect 25872 25162 25924 25168
rect 25884 24954 25912 25162
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25226 24168 25282 24177
rect 25226 24103 25282 24112
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24596 23118 24624 24006
rect 25516 23526 25544 24210
rect 25608 23730 25636 24754
rect 27356 24274 27384 34546
rect 28092 27606 28120 37198
rect 28368 35834 28396 39200
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28552 36718 28580 37198
rect 28540 36712 28592 36718
rect 28540 36654 28592 36660
rect 29092 36712 29144 36718
rect 29092 36654 29144 36660
rect 29104 35834 29132 36654
rect 28356 35828 28408 35834
rect 28356 35770 28408 35776
rect 29092 35828 29144 35834
rect 29092 35770 29144 35776
rect 29276 34672 29328 34678
rect 29276 34614 29328 34620
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 28080 27600 28132 27606
rect 28080 27542 28132 27548
rect 28080 26580 28132 26586
rect 28080 26522 28132 26528
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25700 23866 25728 24074
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 25608 22778 25636 23666
rect 28092 23322 28120 26522
rect 28276 25362 28304 34478
rect 29288 33590 29316 34614
rect 29656 34610 29684 39200
rect 29644 34604 29696 34610
rect 29644 34546 29696 34552
rect 30944 34542 30972 39200
rect 32232 34678 32260 39200
rect 32220 34672 32272 34678
rect 32220 34614 32272 34620
rect 30932 34536 30984 34542
rect 30932 34478 30984 34484
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 32312 28552 32364 28558
rect 32312 28494 32364 28500
rect 32324 28082 32352 28494
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 31772 27470 31800 28018
rect 32876 28014 32904 39200
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35346 37496 35402 37505
rect 35346 37431 35402 37440
rect 36176 37460 36228 37466
rect 35360 37398 35388 37431
rect 36176 37402 36228 37408
rect 35348 37392 35400 37398
rect 35348 37334 35400 37340
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33796 36786 33824 37198
rect 34808 36786 34836 37266
rect 35348 37188 35400 37194
rect 35348 37130 35400 37136
rect 33784 36780 33836 36786
rect 33784 36722 33836 36728
rect 34796 36780 34848 36786
rect 34796 36722 34848 36728
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35360 36378 35388 37130
rect 35348 36372 35400 36378
rect 35348 36314 35400 36320
rect 34888 36168 34940 36174
rect 34888 36110 34940 36116
rect 35440 36168 35492 36174
rect 35440 36110 35492 36116
rect 35624 36168 35676 36174
rect 35624 36110 35676 36116
rect 34900 35698 34928 36110
rect 34888 35692 34940 35698
rect 34888 35634 34940 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 35452 35086 35480 36110
rect 35532 35624 35584 35630
rect 35532 35566 35584 35572
rect 35544 35290 35572 35566
rect 35532 35284 35584 35290
rect 35532 35226 35584 35232
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34888 30728 34940 30734
rect 34888 30670 34940 30676
rect 34900 30258 34928 30670
rect 34888 30252 34940 30258
rect 34888 30194 34940 30200
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 33324 28212 33376 28218
rect 33324 28154 33376 28160
rect 32496 28008 32548 28014
rect 32496 27950 32548 27956
rect 32864 28008 32916 28014
rect 32864 27950 32916 27956
rect 32508 27674 32536 27950
rect 32496 27668 32548 27674
rect 32496 27610 32548 27616
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 33336 25906 33364 28154
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 28264 25356 28316 25362
rect 28264 25298 28316 25304
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 28080 23316 28132 23322
rect 28080 23258 28132 23264
rect 28092 23118 28120 23258
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 28184 22642 28212 23734
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28368 22710 28396 22918
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 30012 22568 30064 22574
rect 30012 22510 30064 22516
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 23216 20602 23244 20742
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23216 19922 23244 20538
rect 23400 20534 23428 21354
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20534 24256 20742
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 24584 19780 24636 19786
rect 24584 19722 24636 19728
rect 22572 19306 22692 19334
rect 22664 6914 22692 19306
rect 22296 6886 22416 6914
rect 22572 6886 22692 6914
rect 22296 3942 22324 6886
rect 22572 4146 22600 6886
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21928 800 21956 3334
rect 23676 3126 23704 3946
rect 23860 3398 23888 19722
rect 24596 19514 24624 19722
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23952 5370 23980 19314
rect 25884 6914 25912 20334
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27264 17746 27292 18022
rect 27632 17814 27660 18022
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27252 17740 27304 17746
rect 27252 17682 27304 17688
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 25608 6886 25912 6914
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 25148 870 25360 898
rect 25148 800 25176 870
rect 3436 734 3740 762
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25332 762 25360 870
rect 25608 762 25636 6886
rect 28920 3738 28948 17546
rect 29552 17128 29604 17134
rect 29552 17070 29604 17076
rect 29564 16794 29592 17070
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 30024 1358 30052 22510
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 31772 20942 31800 21490
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 19854 31800 20878
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 32312 19712 32364 19718
rect 32312 19654 32364 19660
rect 32324 19446 32352 19654
rect 32312 19440 32364 19446
rect 32312 19382 32364 19388
rect 31760 19236 31812 19242
rect 31760 19178 31812 19184
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 30840 3460 30892 3466
rect 30840 3402 30892 3408
rect 30852 3194 30880 3402
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31036 2650 31064 3470
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31312 3058 31340 3402
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 30012 1352 30064 1358
rect 30012 1294 30064 1300
rect 31588 800 31616 3538
rect 25332 734 25636 762
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 31546 0 31658 800
rect 31772 762 31800 19178
rect 31852 4140 31904 4146
rect 31852 4082 31904 4088
rect 31864 3670 31892 4082
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 32588 3936 32640 3942
rect 32588 3878 32640 3884
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 32324 2514 32352 3878
rect 32600 3058 32628 3878
rect 33336 3534 33364 25842
rect 34716 25838 34744 26318
rect 35452 26234 35480 35022
rect 35452 26206 35572 26234
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35544 23322 35572 26206
rect 35532 23316 35584 23322
rect 35532 23258 35584 23264
rect 35636 23254 35664 36110
rect 36188 35154 36216 37402
rect 36740 37262 36768 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 36820 37256 36872 37262
rect 36820 37198 36872 37204
rect 36268 36576 36320 36582
rect 36268 36518 36320 36524
rect 36452 36576 36504 36582
rect 36452 36518 36504 36524
rect 36280 36242 36308 36518
rect 36464 36242 36492 36518
rect 36832 36310 36860 37198
rect 37200 36786 37228 38791
rect 37188 36780 37240 36786
rect 37188 36722 37240 36728
rect 36820 36304 36872 36310
rect 36820 36246 36872 36252
rect 36268 36236 36320 36242
rect 36268 36178 36320 36184
rect 36452 36236 36504 36242
rect 36452 36178 36504 36184
rect 36726 36136 36782 36145
rect 36726 36071 36782 36080
rect 36452 36032 36504 36038
rect 36452 35974 36504 35980
rect 36464 35154 36492 35974
rect 36740 35766 36768 36071
rect 36728 35760 36780 35766
rect 36728 35702 36780 35708
rect 36176 35148 36228 35154
rect 36176 35090 36228 35096
rect 36452 35148 36504 35154
rect 36452 35090 36504 35096
rect 36452 34536 36504 34542
rect 36452 34478 36504 34484
rect 36268 34400 36320 34406
rect 36268 34342 36320 34348
rect 36280 34066 36308 34342
rect 36464 34066 36492 34478
rect 36268 34060 36320 34066
rect 36268 34002 36320 34008
rect 36452 34060 36504 34066
rect 36452 34002 36504 34008
rect 36544 33312 36596 33318
rect 36544 33254 36596 33260
rect 36556 32978 36584 33254
rect 36544 32972 36596 32978
rect 36544 32914 36596 32920
rect 36636 32836 36688 32842
rect 36636 32778 36688 32784
rect 36648 32570 36676 32778
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 36268 32224 36320 32230
rect 36268 32166 36320 32172
rect 36452 32224 36504 32230
rect 36452 32166 36504 32172
rect 36280 31890 36308 32166
rect 36464 31890 36492 32166
rect 36268 31884 36320 31890
rect 36268 31826 36320 31832
rect 36452 31884 36504 31890
rect 36452 31826 36504 31832
rect 36176 31816 36228 31822
rect 36176 31758 36228 31764
rect 35806 31376 35862 31385
rect 35806 31311 35862 31320
rect 35820 31278 35848 31311
rect 36188 31278 36216 31758
rect 35808 31272 35860 31278
rect 35808 31214 35860 31220
rect 36176 31272 36228 31278
rect 36176 31214 36228 31220
rect 37384 30802 37412 39200
rect 37464 37120 37516 37126
rect 37464 37062 37516 37068
rect 37476 36854 37504 37062
rect 37464 36848 37516 36854
rect 37464 36790 37516 36796
rect 38028 35894 38056 39200
rect 38106 36816 38162 36825
rect 38106 36751 38162 36760
rect 38120 36242 38148 36751
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 38028 35866 38148 35894
rect 38016 35692 38068 35698
rect 38016 35634 38068 35640
rect 38028 35465 38056 35634
rect 38014 35456 38070 35465
rect 38014 35391 38070 35400
rect 38120 35154 38148 35866
rect 38108 35148 38160 35154
rect 38108 35090 38160 35096
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 37476 34610 37504 34886
rect 38106 34776 38162 34785
rect 38106 34711 38162 34720
rect 37464 34604 37516 34610
rect 37464 34546 37516 34552
rect 38120 34066 38148 34711
rect 38108 34060 38160 34066
rect 38108 34002 38160 34008
rect 38016 33516 38068 33522
rect 38016 33458 38068 33464
rect 38028 33425 38056 33458
rect 38014 33416 38070 33425
rect 37832 33380 37884 33386
rect 38014 33351 38070 33360
rect 37832 33322 37884 33328
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37372 30796 37424 30802
rect 37372 30738 37424 30744
rect 36726 30696 36782 30705
rect 36726 30631 36782 30640
rect 37372 30660 37424 30666
rect 36740 30326 36768 30631
rect 37372 30602 37424 30608
rect 37384 30326 37412 30602
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 37372 30320 37424 30326
rect 37372 30262 37424 30268
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37186 30016 37242 30025
rect 37186 29951 37242 29960
rect 37200 29714 37228 29951
rect 37188 29708 37240 29714
rect 37188 29650 37240 29656
rect 37292 29170 37320 30194
rect 37476 29730 37504 31282
rect 37384 29702 37504 29730
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 36452 28960 36504 28966
rect 36452 28902 36504 28908
rect 36464 28626 36492 28902
rect 36452 28620 36504 28626
rect 36452 28562 36504 28568
rect 36268 28552 36320 28558
rect 36268 28494 36320 28500
rect 36280 28082 36308 28494
rect 37384 28098 37412 29702
rect 37464 29572 37516 29578
rect 37464 29514 37516 29520
rect 37476 29306 37504 29514
rect 37464 29300 37516 29306
rect 37464 29242 37516 29248
rect 37464 29164 37516 29170
rect 37464 29106 37516 29112
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 37292 28070 37412 28098
rect 37292 26926 37320 28070
rect 37280 26920 37332 26926
rect 37280 26862 37332 26868
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 35806 25936 35862 25945
rect 36280 25906 36308 26318
rect 37292 25906 37320 26862
rect 37372 26308 37424 26314
rect 37372 26250 37424 26256
rect 37384 26042 37412 26250
rect 37372 26036 37424 26042
rect 37372 25978 37424 25984
rect 35806 25871 35862 25880
rect 36268 25900 36320 25906
rect 35820 25838 35848 25871
rect 36268 25842 36320 25848
rect 37280 25900 37332 25906
rect 37280 25842 37332 25848
rect 35808 25832 35860 25838
rect 35808 25774 35860 25780
rect 37476 25770 37504 29106
rect 37556 29096 37608 29102
rect 37556 29038 37608 29044
rect 37464 25764 37516 25770
rect 37464 25706 37516 25712
rect 36176 25220 36228 25226
rect 36176 25162 36228 25168
rect 35624 23248 35676 23254
rect 35624 23190 35676 23196
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34518 21856 34574 21865
rect 34518 21791 34574 21800
rect 34532 20874 34560 21791
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34520 20868 34572 20874
rect 34520 20810 34572 20816
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35624 19780 35676 19786
rect 35624 19722 35676 19728
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35636 18465 35664 19722
rect 35622 18456 35678 18465
rect 35622 18391 35678 18400
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34520 17128 34572 17134
rect 34518 17096 34520 17105
rect 34572 17096 34574 17105
rect 34518 17031 34574 17040
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34518 14376 34574 14385
rect 34518 14311 34520 14320
rect 34572 14311 34574 14320
rect 34520 14282 34572 14288
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35808 12232 35860 12238
rect 35808 12174 35860 12180
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35820 11354 35848 12174
rect 35808 11348 35860 11354
rect 35808 11290 35860 11296
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 36188 6914 36216 25162
rect 37186 23896 37242 23905
rect 37186 23831 37242 23840
rect 37200 23186 37228 23831
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37292 23254 37320 23666
rect 37280 23248 37332 23254
rect 37280 23190 37332 23196
rect 37188 23180 37240 23186
rect 37188 23122 37240 23128
rect 37476 22794 37504 25706
rect 37568 24857 37596 29038
rect 37554 24848 37610 24857
rect 37554 24783 37610 24792
rect 37384 22766 37504 22794
rect 36544 22432 36596 22438
rect 36544 22374 36596 22380
rect 36636 22432 36688 22438
rect 36636 22374 36688 22380
rect 36556 22098 36584 22374
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 36648 21962 36676 22374
rect 36636 21956 36688 21962
rect 36636 21898 36688 21904
rect 36268 21344 36320 21350
rect 36268 21286 36320 21292
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 36280 21010 36308 21286
rect 36648 21010 36676 21286
rect 36268 21004 36320 21010
rect 36268 20946 36320 20952
rect 36636 21004 36688 21010
rect 36636 20946 36688 20952
rect 37186 20496 37242 20505
rect 37186 20431 37242 20440
rect 37200 19922 37228 20431
rect 37188 19916 37240 19922
rect 37188 19858 37240 19864
rect 37186 15056 37242 15065
rect 37186 14991 37242 15000
rect 37200 14482 37228 14991
rect 37188 14476 37240 14482
rect 37188 14418 37240 14424
rect 37186 13696 37242 13705
rect 37186 13631 37242 13640
rect 37200 13394 37228 13631
rect 37188 13388 37240 13394
rect 37188 13330 37240 13336
rect 37188 12300 37240 12306
rect 37188 12242 37240 12248
rect 36268 11552 36320 11558
rect 36268 11494 36320 11500
rect 36280 11218 36308 11494
rect 36268 11212 36320 11218
rect 36268 11154 36320 11160
rect 37200 10985 37228 12242
rect 37280 12164 37332 12170
rect 37280 12106 37332 12112
rect 37186 10976 37242 10985
rect 37186 10911 37242 10920
rect 37292 10810 37320 12106
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 36268 10464 36320 10470
rect 36268 10406 36320 10412
rect 36280 10130 36308 10406
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 36452 9988 36504 9994
rect 36452 9930 36504 9936
rect 36464 9722 36492 9930
rect 36452 9716 36504 9722
rect 36452 9658 36504 9664
rect 37186 9616 37242 9625
rect 37384 9586 37412 22766
rect 37568 22522 37596 24783
rect 37476 22494 37596 22522
rect 37476 12850 37504 22494
rect 37660 21554 37688 32370
rect 37844 25430 37872 33322
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 38120 32745 38148 32778
rect 38106 32736 38162 32745
rect 38106 32671 38162 32680
rect 37924 32360 37976 32366
rect 37924 32302 37976 32308
rect 37936 30258 37964 32302
rect 38106 32056 38162 32065
rect 38106 31991 38162 32000
rect 38120 31890 38148 31991
rect 38108 31884 38160 31890
rect 38108 31826 38160 31832
rect 38108 31136 38160 31142
rect 38108 31078 38160 31084
rect 37924 30252 37976 30258
rect 37924 30194 37976 30200
rect 37936 25906 37964 30194
rect 38120 29714 38148 31078
rect 38108 29708 38160 29714
rect 38108 29650 38160 29656
rect 38106 29336 38162 29345
rect 38106 29271 38162 29280
rect 38120 28626 38148 29271
rect 38108 28620 38160 28626
rect 38108 28562 38160 28568
rect 38016 26988 38068 26994
rect 38016 26930 38068 26936
rect 38028 26625 38056 26930
rect 38014 26616 38070 26625
rect 38014 26551 38070 26560
rect 38200 26308 38252 26314
rect 38200 26250 38252 26256
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 37924 25696 37976 25702
rect 37924 25638 37976 25644
rect 37832 25424 37884 25430
rect 37832 25366 37884 25372
rect 37936 25362 37964 25638
rect 37924 25356 37976 25362
rect 37924 25298 37976 25304
rect 38108 25288 38160 25294
rect 38108 25230 38160 25236
rect 38120 24818 38148 25230
rect 38108 24812 38160 24818
rect 38108 24754 38160 24760
rect 38108 24200 38160 24206
rect 38108 24142 38160 24148
rect 37924 23520 37976 23526
rect 37924 23462 37976 23468
rect 37936 23186 37964 23462
rect 38120 23186 38148 24142
rect 37924 23180 37976 23186
rect 37924 23122 37976 23128
rect 38108 23180 38160 23186
rect 38108 23122 38160 23128
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37648 16652 37700 16658
rect 37648 16594 37700 16600
rect 37556 16516 37608 16522
rect 37556 16458 37608 16464
rect 37568 16250 37596 16458
rect 37660 16425 37688 16594
rect 37646 16416 37702 16425
rect 37646 16351 37702 16360
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 37568 12986 37596 13194
rect 37556 12980 37608 12986
rect 37556 12922 37608 12928
rect 37660 12866 37688 14962
rect 37752 13002 37780 22578
rect 38106 22536 38162 22545
rect 38106 22471 38162 22480
rect 38120 22098 38148 22471
rect 38108 22092 38160 22098
rect 38108 22034 38160 22040
rect 38106 21176 38162 21185
rect 38106 21111 38162 21120
rect 38120 21010 38148 21111
rect 38108 21004 38160 21010
rect 38108 20946 38160 20952
rect 37924 20256 37976 20262
rect 37924 20198 37976 20204
rect 37936 19922 37964 20198
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38108 19848 38160 19854
rect 38108 19790 38160 19796
rect 38120 19378 38148 19790
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38120 16658 38148 16934
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 38108 15496 38160 15502
rect 38108 15438 38160 15444
rect 37924 14816 37976 14822
rect 37924 14758 37976 14764
rect 37936 14482 37964 14758
rect 38120 14482 38148 15438
rect 37924 14476 37976 14482
rect 37924 14418 37976 14424
rect 38108 14476 38160 14482
rect 38108 14418 38160 14424
rect 37832 13728 37884 13734
rect 37832 13670 37884 13676
rect 37844 13394 37872 13670
rect 37832 13388 37884 13394
rect 37832 13330 37884 13336
rect 37752 12974 37872 13002
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37568 12838 37688 12866
rect 37740 12844 37792 12850
rect 37186 9551 37242 9560
rect 37372 9580 37424 9586
rect 37200 9042 37228 9551
rect 37372 9522 37424 9528
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37568 6914 37596 12838
rect 37740 12786 37792 12792
rect 37648 11552 37700 11558
rect 37648 11494 37700 11500
rect 37660 11218 37688 11494
rect 37648 11212 37700 11218
rect 37648 11154 37700 11160
rect 36188 6886 36308 6914
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 36280 5545 36308 6886
rect 37292 6886 37596 6914
rect 36266 5536 36322 5545
rect 36266 5471 36322 5480
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 37188 4684 37240 4690
rect 37188 4626 37240 4632
rect 37200 4185 37228 4626
rect 37186 4176 37242 4185
rect 37292 4146 37320 6886
rect 37186 4111 37242 4120
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37752 4078 37780 12786
rect 37844 11762 37872 12974
rect 37832 11756 37884 11762
rect 37832 11698 37884 11704
rect 37844 11082 37872 11698
rect 38106 11656 38162 11665
rect 38106 11591 38162 11600
rect 38120 11218 38148 11591
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 37832 11076 37884 11082
rect 37832 11018 37884 11024
rect 37844 10674 37872 11018
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38120 10130 38148 10231
rect 38108 10124 38160 10130
rect 38108 10066 38160 10072
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 37936 9042 37964 9318
rect 37924 9036 37976 9042
rect 37924 8978 37976 8984
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8498 38148 8910
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38108 5024 38160 5030
rect 38108 4966 38160 4972
rect 38120 4690 38148 4966
rect 38108 4684 38160 4690
rect 38108 4626 38160 4632
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37936 4282 37964 4490
rect 37924 4276 37976 4282
rect 37924 4218 37976 4224
rect 34520 4072 34572 4078
rect 34520 4014 34572 4020
rect 37740 4072 37792 4078
rect 37740 4014 37792 4020
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 32784 3126 32812 3334
rect 32772 3120 32824 3126
rect 32772 3062 32824 3068
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 33336 2990 33364 3470
rect 34152 3460 34204 3466
rect 34152 3402 34204 3408
rect 33324 2984 33376 2990
rect 33324 2926 33376 2932
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32496 2848 32548 2854
rect 32496 2790 32548 2796
rect 32508 2514 32536 2790
rect 32312 2508 32364 2514
rect 32312 2450 32364 2456
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 32864 2508 32916 2514
rect 32864 2450 32916 2456
rect 32048 870 32260 898
rect 32048 762 32076 870
rect 32232 800 32260 870
rect 32876 800 32904 2450
rect 33520 800 33548 2926
rect 34164 800 34192 3402
rect 34532 2145 34560 4014
rect 35716 4004 35768 4010
rect 35716 3946 35768 3952
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 35624 3936 35676 3942
rect 35624 3878 35676 3884
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 2378 34652 3334
rect 34716 2514 34744 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35360 3126 35388 3878
rect 35636 3194 35664 3878
rect 35728 3194 35756 3946
rect 37832 3936 37884 3942
rect 37832 3878 37884 3884
rect 37372 3664 37424 3670
rect 37372 3606 37424 3612
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 35716 3188 35768 3194
rect 35716 3130 35768 3136
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34704 2508 34756 2514
rect 34704 2450 34756 2456
rect 34612 2372 34664 2378
rect 34612 2314 34664 2320
rect 34518 2136 34574 2145
rect 34518 2071 34574 2080
rect 34520 1352 34572 1358
rect 34520 1294 34572 1300
rect 31772 734 32076 762
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34532 785 34560 1294
rect 35452 800 35480 2926
rect 36832 1714 36860 3538
rect 37188 2372 37240 2378
rect 37188 2314 37240 2320
rect 36740 1686 36860 1714
rect 36740 800 36768 1686
rect 34518 776 34574 785
rect 34518 711 34574 720
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 37200 105 37228 2314
rect 37384 800 37412 3606
rect 37844 3602 37872 3878
rect 37832 3596 37884 3602
rect 37832 3538 37884 3544
rect 38014 3496 38070 3505
rect 37464 3460 37516 3466
rect 38014 3431 38070 3440
rect 37464 3402 37516 3408
rect 37476 2650 37504 3402
rect 38028 3126 38056 3431
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38212 2972 38240 26250
rect 38660 3392 38712 3398
rect 38660 3334 38712 3340
rect 38028 2944 38240 2972
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38028 800 38056 2944
rect 38672 800 38700 3334
rect 37186 96 37242 105
rect 37186 31 37242 40
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
<< via2 >>
rect 3330 38800 3386 38856
rect 1398 36760 1454 36816
rect 1858 32000 1914 32056
rect 2778 34720 2834 34776
rect 1858 23160 1914 23216
rect 3422 37460 3478 37496
rect 3422 37440 3424 37460
rect 3424 37440 3476 37460
rect 3476 37440 3478 37460
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 3698 36080 3754 36136
rect 3422 33360 3478 33416
rect 3514 25880 3570 25936
rect 1858 19760 1914 19816
rect 2134 19080 2190 19136
rect 1582 15680 1638 15736
rect 1398 15000 1454 15056
rect 1398 14356 1400 14376
rect 1400 14356 1452 14376
rect 1452 14356 1454 14376
rect 1398 14320 1454 14356
rect 1858 13640 1914 13696
rect 1858 8880 1914 8936
rect 1398 7520 1454 7576
rect 2042 6196 2044 6216
rect 2044 6196 2096 6216
rect 2096 6196 2098 6216
rect 2042 6160 2098 6196
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 3330 4120 3386 4176
rect 2778 2760 2834 2816
rect 2870 2080 2926 2136
rect 3330 1400 3386 1456
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3514 4800 3570 4856
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8200 4122 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3514 3440 3570 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 18418 24112 18474 24168
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 18786 24248 18842 24304
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20534 24812 20590 24848
rect 20534 24792 20536 24812
rect 20536 24792 20588 24812
rect 20588 24792 20590 24812
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24674 24248 24730 24304
rect 25226 24112 25282 24168
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35346 37440 35402 37496
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 37186 38800 37242 38856
rect 36726 36080 36782 36136
rect 35806 31320 35862 31376
rect 38106 36760 38162 36816
rect 38014 35400 38070 35456
rect 38106 34720 38162 34776
rect 38014 33360 38070 33416
rect 36726 30640 36782 30696
rect 37186 29960 37242 30016
rect 35806 25880 35862 25936
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34518 21800 34574 21856
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35622 18400 35678 18456
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34518 17076 34520 17096
rect 34520 17076 34572 17096
rect 34572 17076 34574 17096
rect 34518 17040 34574 17076
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34518 14340 34574 14376
rect 34518 14320 34520 14340
rect 34520 14320 34572 14340
rect 34572 14320 34574 14340
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37186 23840 37242 23896
rect 37554 24792 37610 24848
rect 37186 20440 37242 20496
rect 37186 15000 37242 15056
rect 37186 13640 37242 13696
rect 37186 10920 37242 10976
rect 37186 9560 37242 9616
rect 38106 32680 38162 32736
rect 38106 32000 38162 32056
rect 38106 29280 38162 29336
rect 38014 26560 38070 26616
rect 37646 16360 37702 16416
rect 38106 22480 38162 22536
rect 38106 21120 38162 21176
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 36266 5480 36322 5536
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37186 4120 37242 4176
rect 38106 11600 38162 11656
rect 38106 10240 38162 10296
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 34518 2080 34574 2136
rect 34518 720 34574 776
rect 38014 3440 38070 3496
rect 37186 40 37242 96
<< metal3 >>
rect 0 39388 800 39628
rect 0 38858 800 38948
rect 3325 38858 3391 38861
rect 0 38856 3391 38858
rect 0 38800 3330 38856
rect 3386 38800 3391 38856
rect 0 38798 3391 38800
rect 0 38708 800 38798
rect 3325 38795 3391 38798
rect 37181 38858 37247 38861
rect 39200 38858 40000 38948
rect 37181 38856 40000 38858
rect 37181 38800 37186 38856
rect 37242 38800 40000 38856
rect 37181 38798 40000 38800
rect 37181 38795 37247 38798
rect 39200 38708 40000 38798
rect 39200 38028 40000 38268
rect 0 37498 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 3417 37498 3483 37501
rect 0 37496 3483 37498
rect 0 37440 3422 37496
rect 3478 37440 3483 37496
rect 0 37438 3483 37440
rect 0 37348 800 37438
rect 3417 37435 3483 37438
rect 35341 37498 35407 37501
rect 39200 37498 40000 37588
rect 35341 37496 40000 37498
rect 35341 37440 35346 37496
rect 35402 37440 40000 37496
rect 35341 37438 40000 37440
rect 35341 37435 35407 37438
rect 39200 37348 40000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 1393 36818 1459 36821
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 0 36668 800 36758
rect 1393 36755 1459 36758
rect 38101 36818 38167 36821
rect 39200 36818 40000 36908
rect 38101 36816 40000 36818
rect 38101 36760 38106 36816
rect 38162 36760 40000 36816
rect 38101 36758 40000 36760
rect 38101 36755 38167 36758
rect 39200 36668 40000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36228
rect 3693 36138 3759 36141
rect 0 36136 3759 36138
rect 0 36080 3698 36136
rect 3754 36080 3759 36136
rect 0 36078 3759 36080
rect 0 35988 800 36078
rect 3693 36075 3759 36078
rect 36721 36138 36787 36141
rect 39200 36138 40000 36228
rect 36721 36136 40000 36138
rect 36721 36080 36726 36136
rect 36782 36080 40000 36136
rect 36721 36078 40000 36080
rect 36721 36075 36787 36078
rect 39200 35988 40000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35308 800 35548
rect 38009 35458 38075 35461
rect 39200 35458 40000 35548
rect 38009 35456 40000 35458
rect 38009 35400 38014 35456
rect 38070 35400 40000 35456
rect 38009 35398 40000 35400
rect 38009 35395 38075 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 39200 35308 40000 35398
rect 0 34778 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 2773 34778 2839 34781
rect 0 34776 2839 34778
rect 0 34720 2778 34776
rect 2834 34720 2839 34776
rect 0 34718 2839 34720
rect 0 34628 800 34718
rect 2773 34715 2839 34718
rect 38101 34778 38167 34781
rect 39200 34778 40000 34868
rect 38101 34776 40000 34778
rect 38101 34720 38106 34776
rect 38162 34720 40000 34776
rect 38101 34718 40000 34720
rect 38101 34715 38167 34718
rect 39200 34628 40000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 3417 33418 3483 33421
rect 0 33416 3483 33418
rect 0 33360 3422 33416
rect 3478 33360 3483 33416
rect 0 33358 3483 33360
rect 0 33268 800 33358
rect 3417 33355 3483 33358
rect 38009 33418 38075 33421
rect 39200 33418 40000 33508
rect 38009 33416 40000 33418
rect 38009 33360 38014 33416
rect 38070 33360 40000 33416
rect 38009 33358 40000 33360
rect 38009 33355 38075 33358
rect 39200 33268 40000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 38101 32738 38167 32741
rect 39200 32738 40000 32828
rect 38101 32736 40000 32738
rect 38101 32680 38106 32736
rect 38162 32680 40000 32736
rect 38101 32678 40000 32680
rect 38101 32675 38167 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 39200 32588 40000 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 38101 32058 38167 32061
rect 39200 32058 40000 32148
rect 38101 32056 40000 32058
rect 38101 32000 38106 32056
rect 38162 32000 40000 32056
rect 38101 31998 40000 32000
rect 38101 31995 38167 31998
rect 39200 31908 40000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31228 800 31468
rect 35801 31378 35867 31381
rect 39200 31378 40000 31468
rect 35801 31376 40000 31378
rect 35801 31320 35806 31376
rect 35862 31320 40000 31376
rect 35801 31318 40000 31320
rect 35801 31315 35867 31318
rect 39200 31228 40000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 36721 30698 36787 30701
rect 39200 30698 40000 30788
rect 36721 30696 40000 30698
rect 36721 30640 36726 30696
rect 36782 30640 40000 30696
rect 36721 30638 40000 30640
rect 36721 30635 36787 30638
rect 39200 30548 40000 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 37181 30018 37247 30021
rect 39200 30018 40000 30108
rect 37181 30016 40000 30018
rect 37181 29960 37186 30016
rect 37242 29960 40000 30016
rect 37181 29958 40000 29960
rect 37181 29955 37247 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 39200 29868 40000 29958
rect 0 29188 800 29428
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 38101 29338 38167 29341
rect 39200 29338 40000 29428
rect 38101 29336 40000 29338
rect 38101 29280 38106 29336
rect 38162 29280 40000 29336
rect 38101 29278 40000 29280
rect 38101 29275 38167 29278
rect 39200 29188 40000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28508 800 28748
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 39200 27828 40000 28068
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 39200 27148 40000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 38009 26618 38075 26621
rect 39200 26618 40000 26708
rect 38009 26616 40000 26618
rect 38009 26560 38014 26616
rect 38070 26560 40000 26616
rect 38009 26558 40000 26560
rect 38009 26555 38075 26558
rect 39200 26468 40000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 26028
rect 3509 25938 3575 25941
rect 0 25936 3575 25938
rect 0 25880 3514 25936
rect 3570 25880 3575 25936
rect 0 25878 3575 25880
rect 0 25788 800 25878
rect 3509 25875 3575 25878
rect 35801 25938 35867 25941
rect 39200 25938 40000 26028
rect 35801 25936 40000 25938
rect 35801 25880 35806 25936
rect 35862 25880 40000 25936
rect 35801 25878 40000 25880
rect 35801 25875 35867 25878
rect 39200 25788 40000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25108 800 25348
rect 39200 25108 40000 25348
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 20529 24850 20595 24853
rect 37549 24850 37615 24853
rect 20529 24848 37615 24850
rect 20529 24792 20534 24848
rect 20590 24792 37554 24848
rect 37610 24792 37615 24848
rect 20529 24790 37615 24792
rect 20529 24787 20595 24790
rect 37549 24787 37615 24790
rect 0 24428 800 24668
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 39200 24428 40000 24668
rect 18781 24306 18847 24309
rect 24669 24306 24735 24309
rect 18781 24304 24735 24306
rect 18781 24248 18786 24304
rect 18842 24248 24674 24304
rect 24730 24248 24735 24304
rect 18781 24246 24735 24248
rect 18781 24243 18847 24246
rect 24669 24243 24735 24246
rect 18413 24170 18479 24173
rect 25221 24170 25287 24173
rect 18413 24168 25287 24170
rect 18413 24112 18418 24168
rect 18474 24112 25226 24168
rect 25282 24112 25287 24168
rect 18413 24110 25287 24112
rect 18413 24107 18479 24110
rect 25221 24107 25287 24110
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 37181 23898 37247 23901
rect 39200 23898 40000 23988
rect 37181 23896 40000 23898
rect 37181 23840 37186 23896
rect 37242 23840 40000 23896
rect 37181 23838 40000 23840
rect 37181 23835 37247 23838
rect 39200 23748 40000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 38101 22538 38167 22541
rect 39200 22538 40000 22628
rect 38101 22536 40000 22538
rect 38101 22480 38106 22536
rect 38162 22480 40000 22536
rect 38101 22478 40000 22480
rect 38101 22475 38167 22478
rect 39200 22388 40000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 34513 21858 34579 21861
rect 39200 21858 40000 21948
rect 34513 21856 40000 21858
rect 34513 21800 34518 21856
rect 34574 21800 40000 21856
rect 34513 21798 40000 21800
rect 34513 21795 34579 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 39200 21708 40000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 38101 21178 38167 21181
rect 39200 21178 40000 21268
rect 38101 21176 40000 21178
rect 38101 21120 38106 21176
rect 38162 21120 40000 21176
rect 38101 21118 40000 21120
rect 38101 21115 38167 21118
rect 39200 21028 40000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 37181 20498 37247 20501
rect 39200 20498 40000 20588
rect 37181 20496 40000 20498
rect 37181 20440 37186 20496
rect 37242 20440 40000 20496
rect 37181 20438 40000 20440
rect 37181 20435 37247 20438
rect 39200 20348 40000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19668 800 19758
rect 1853 19755 1919 19758
rect 39200 19668 40000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2129 19138 2195 19141
rect 0 19136 2195 19138
rect 0 19080 2134 19136
rect 2190 19080 2195 19136
rect 0 19078 2195 19080
rect 0 18988 800 19078
rect 2129 19075 2195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 39200 18988 40000 19228
rect 0 18308 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 35617 18458 35683 18461
rect 39200 18458 40000 18548
rect 35617 18456 40000 18458
rect 35617 18400 35622 18456
rect 35678 18400 40000 18456
rect 35617 18398 40000 18400
rect 35617 18395 35683 18398
rect 39200 18308 40000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17628 800 17718
rect 2773 17715 2839 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 16948 800 17188
rect 34513 17098 34579 17101
rect 39200 17098 40000 17188
rect 34513 17096 40000 17098
rect 34513 17040 34518 17096
rect 34574 17040 40000 17096
rect 34513 17038 40000 17040
rect 34513 17035 34579 17038
rect 39200 16948 40000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 37641 16418 37707 16421
rect 39200 16418 40000 16508
rect 37641 16416 40000 16418
rect 37641 16360 37646 16416
rect 37702 16360 40000 16416
rect 37641 16358 40000 16360
rect 37641 16355 37707 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 39200 16268 40000 16358
rect 0 15738 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 1577 15738 1643 15741
rect 0 15736 1643 15738
rect 0 15680 1582 15736
rect 1638 15680 1643 15736
rect 0 15678 1643 15680
rect 0 15588 800 15678
rect 1577 15675 1643 15678
rect 39200 15588 40000 15828
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14908 800 14998
rect 1393 14995 1459 14998
rect 37181 15058 37247 15061
rect 39200 15058 40000 15148
rect 37181 15056 40000 15058
rect 37181 15000 37186 15056
rect 37242 15000 40000 15056
rect 37181 14998 40000 15000
rect 37181 14995 37247 14998
rect 39200 14908 40000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14378 800 14468
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14228 800 14318
rect 1393 14315 1459 14318
rect 34513 14378 34579 14381
rect 39200 14378 40000 14468
rect 34513 14376 40000 14378
rect 34513 14320 34518 14376
rect 34574 14320 40000 14376
rect 34513 14318 40000 14320
rect 34513 14315 34579 14318
rect 39200 14228 40000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 1853 13698 1919 13701
rect 0 13696 1919 13698
rect 0 13640 1858 13696
rect 1914 13640 1919 13696
rect 0 13638 1919 13640
rect 0 13548 800 13638
rect 1853 13635 1919 13638
rect 37181 13698 37247 13701
rect 39200 13698 40000 13788
rect 37181 13696 40000 13698
rect 37181 13640 37186 13696
rect 37242 13640 40000 13696
rect 37181 13638 40000 13640
rect 37181 13635 37247 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 39200 13548 40000 13638
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 39200 12868 40000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12188 800 12278
rect 2773 12275 2839 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11658 800 11748
rect 2773 11658 2839 11661
rect 0 11656 2839 11658
rect 0 11600 2778 11656
rect 2834 11600 2839 11656
rect 0 11598 2839 11600
rect 0 11508 800 11598
rect 2773 11595 2839 11598
rect 38101 11658 38167 11661
rect 39200 11658 40000 11748
rect 38101 11656 40000 11658
rect 38101 11600 38106 11656
rect 38162 11600 40000 11656
rect 38101 11598 40000 11600
rect 38101 11595 38167 11598
rect 39200 11508 40000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 37181 10978 37247 10981
rect 39200 10978 40000 11068
rect 37181 10976 40000 10978
rect 37181 10920 37186 10976
rect 37242 10920 40000 10976
rect 37181 10918 40000 10920
rect 37181 10915 37247 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 39200 10828 40000 10918
rect 0 10148 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 38101 10298 38167 10301
rect 39200 10298 40000 10388
rect 38101 10296 40000 10298
rect 38101 10240 38106 10296
rect 38162 10240 40000 10296
rect 38101 10238 40000 10240
rect 38101 10235 38167 10238
rect 39200 10148 40000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 37181 9618 37247 9621
rect 39200 9618 40000 9708
rect 37181 9616 40000 9618
rect 37181 9560 37186 9616
rect 37242 9560 40000 9616
rect 37181 9558 40000 9560
rect 37181 9555 37247 9558
rect 39200 9468 40000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 9028
rect 1853 8938 1919 8941
rect 0 8936 1919 8938
rect 0 8880 1858 8936
rect 1914 8880 1919 8936
rect 0 8878 1919 8880
rect 0 8788 800 8878
rect 1853 8875 1919 8878
rect 39200 8788 40000 9028
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8348
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8108 800 8198
rect 4061 8195 4127 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 39200 8108 40000 8348
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7428 800 7518
rect 1393 7515 1459 7518
rect 39200 7428 40000 7668
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6748 800 6988
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6308
rect 2037 6218 2103 6221
rect 0 6216 2103 6218
rect 0 6160 2042 6216
rect 2098 6160 2103 6216
rect 0 6158 2103 6160
rect 0 6068 800 6158
rect 2037 6155 2103 6158
rect 39200 6068 40000 6308
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 36261 5538 36327 5541
rect 39200 5538 40000 5628
rect 36261 5536 40000 5538
rect 36261 5480 36266 5536
rect 36322 5480 40000 5536
rect 36261 5478 40000 5480
rect 36261 5475 36327 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 39200 5388 40000 5478
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 3509 4858 3575 4861
rect 0 4856 3575 4858
rect 0 4800 3514 4856
rect 3570 4800 3575 4856
rect 0 4798 3575 4800
rect 0 4708 800 4798
rect 3509 4795 3575 4798
rect 39200 4708 40000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4268
rect 3325 4178 3391 4181
rect 0 4176 3391 4178
rect 0 4120 3330 4176
rect 3386 4120 3391 4176
rect 0 4118 3391 4120
rect 0 4028 800 4118
rect 3325 4115 3391 4118
rect 37181 4178 37247 4181
rect 39200 4178 40000 4268
rect 37181 4176 40000 4178
rect 37181 4120 37186 4176
rect 37242 4120 40000 4176
rect 37181 4118 40000 4120
rect 37181 4115 37247 4118
rect 39200 4028 40000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 3509 3498 3575 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 0 3348 800 3438
rect 3509 3435 3575 3438
rect 38009 3498 38075 3501
rect 39200 3498 40000 3588
rect 38009 3496 40000 3498
rect 38009 3440 38014 3496
rect 38070 3440 40000 3496
rect 38009 3438 40000 3440
rect 38009 3435 38075 3438
rect 39200 3348 40000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2818 800 2908
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2668 800 2758
rect 2773 2755 2839 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 39200 2668 40000 2908
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 1988 800 2078
rect 2865 2075 2931 2078
rect 34513 2138 34579 2141
rect 39200 2138 40000 2228
rect 34513 2136 40000 2138
rect 34513 2080 34518 2136
rect 34574 2080 40000 2136
rect 34513 2078 40000 2080
rect 34513 2075 34579 2078
rect 39200 1988 40000 2078
rect 0 1458 800 1548
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1308 800 1398
rect 3325 1395 3391 1398
rect 0 628 800 868
rect 34513 778 34579 781
rect 39200 778 40000 868
rect 34513 776 40000 778
rect 34513 720 34518 776
rect 34574 720 40000 776
rect 34513 718 40000 720
rect 34513 715 34579 718
rect 39200 628 40000 718
rect 37181 98 37247 101
rect 39200 98 40000 188
rect 37181 96 40000 98
rect 37181 40 37186 96
rect 37242 40 40000 96
rect 37181 38 40000 40
rect 37181 35 37247 38
rect 39200 -52 40000 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1644511149
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_147
timestamp 1644511149
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_179
timestamp 1644511149
transform 1 0 17572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1644511149
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_228
timestamp 1644511149
transform 1 0 22080 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1644511149
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_396
timestamp 1644511149
transform 1 0 37536 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1644511149
transform 1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1644511149
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_246
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_258
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_270
timestamp 1644511149
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1644511149
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_321
timestamp 1644511149
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_341
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1644511149
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_120
timestamp 1644511149
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_147
timestamp 1644511149
transform 1 0 14628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1644511149
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1644511149
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_375
timestamp 1644511149
transform 1 0 35604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_402
timestamp 1644511149
transform 1 0 38088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_202
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_240
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1644511149
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_355
timestamp 1644511149
transform 1 0 33764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_359
timestamp 1644511149
transform 1 0 34132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_371
timestamp 1644511149
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_378
timestamp 1644511149
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_382
timestamp 1644511149
transform 1 0 36248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1644511149
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_398
timestamp 1644511149
transform 1 0 37720 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1644511149
transform 1 0 38456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_8
timestamp 1644511149
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1644511149
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_122
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1644511149
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1644511149
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_202
timestamp 1644511149
transform 1 0 19688 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_210
timestamp 1644511149
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_216
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_228
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_381
timestamp 1644511149
transform 1 0 36156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1644511149
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1644511149
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_400
timestamp 1644511149
transform 1 0 37904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_11
timestamp 1644511149
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_8
timestamp 1644511149
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1644511149
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1644511149
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1644511149
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1644511149
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_88
timestamp 1644511149
transform 1 0 9200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_100
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_112
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_124
timestamp 1644511149
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_231
timestamp 1644511149
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1644511149
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1644511149
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_95
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1644511149
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1644511149
transform 1 0 37904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1644511149
transform 1 0 38456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_8
timestamp 1644511149
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_20
timestamp 1644511149
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1644511149
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1644511149
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_397
timestamp 1644511149
transform 1 0 37628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1644511149
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_73
timestamp 1644511149
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1644511149
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_381
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_9
timestamp 1644511149
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_21
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_33
timestamp 1644511149
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1644511149
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1644511149
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_60
timestamp 1644511149
transform 1 0 6624 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_72
timestamp 1644511149
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_84
timestamp 1644511149
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_96
timestamp 1644511149
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1644511149
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_398
timestamp 1644511149
transform 1 0 37720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_406
timestamp 1644511149
transform 1 0 38456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_12
timestamp 1644511149
transform 1 0 2208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_210
timestamp 1644511149
transform 1 0 20424 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_222
timestamp 1644511149
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_234
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_373
timestamp 1644511149
transform 1 0 35420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_378
timestamp 1644511149
transform 1 0 35880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1644511149
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_399
timestamp 1644511149
transform 1 0 37812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 1644511149
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_18
timestamp 1644511149
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1644511149
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1644511149
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1644511149
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1644511149
transform 1 0 38456 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_8
timestamp 1644511149
transform 1 0 1840 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1644511149
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1644511149
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_381
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_29
timestamp 1644511149
transform 1 0 3772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_41
timestamp 1644511149
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_400
timestamp 1644511149
transform 1 0 37904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1644511149
transform 1 0 38456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1644511149
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_224
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_236
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_37
timestamp 1644511149
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1644511149
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_206
timestamp 1644511149
transform 1 0 20056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1644511149
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_398
timestamp 1644511149
transform 1 0 37720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1644511149
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_400
timestamp 1644511149
transform 1 0 37904 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1644511149
transform 1 0 38456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1644511149
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1644511149
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1644511149
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1644511149
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1644511149
transform 1 0 29808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_348
timestamp 1644511149
transform 1 0 33120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1644511149
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1644511149
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_400
timestamp 1644511149
transform 1 0 37904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1644511149
transform 1 0 38456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1644511149
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_8
timestamp 1644511149
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1644511149
transform 1 0 22448 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_244
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_268
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_284
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_291
timestamp 1644511149
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_315
timestamp 1644511149
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1644511149
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_9
timestamp 1644511149
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1644511149
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1644511149
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1644511149
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_358
timestamp 1644511149
transform 1 0 34040 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_370
timestamp 1644511149
transform 1 0 35144 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_382
timestamp 1644511149
transform 1 0 36248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1644511149
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1644511149
transform 1 0 37904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1644511149
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_217
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_274
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_336
timestamp 1644511149
transform 1 0 32016 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_348
timestamp 1644511149
transform 1 0 33120 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1644511149
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 1644511149
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1644511149
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1644511149
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1644511149
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1644511149
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_243
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1644511149
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_398
timestamp 1644511149
transform 1 0 37720 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1644511149
transform 1 0 38456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1644511149
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_256
timestamp 1644511149
transform 1 0 24656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_268
timestamp 1644511149
transform 1 0 25760 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_381
timestamp 1644511149
transform 1 0 36156 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_201
timestamp 1644511149
transform 1 0 19596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_232
timestamp 1644511149
transform 1 0 22448 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_243
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_255
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_267
timestamp 1644511149
transform 1 0 25668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_398
timestamp 1644511149
transform 1 0 37720 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1644511149
transform 1 0 38456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_210
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_222
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_234
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1644511149
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_381
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1644511149
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_228
timestamp 1644511149
transform 1 0 22080 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_235
timestamp 1644511149
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_247
timestamp 1644511149
transform 1 0 23828 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_315
timestamp 1644511149
transform 1 0 30084 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_399
timestamp 1644511149
transform 1 0 37812 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1644511149
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1644511149
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1644511149
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_293
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_297
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1644511149
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1644511149
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1644511149
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1644511149
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_244
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_256
timestamp 1644511149
transform 1 0 24656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1644511149
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1644511149
transform 1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_12
timestamp 1644511149
transform 1 0 2208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1644511149
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_211
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_236
timestamp 1644511149
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_286
timestamp 1644511149
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_298
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1644511149
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_400
timestamp 1644511149
transform 1 0 37904 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1644511149
transform 1 0 38456 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_198
timestamp 1644511149
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_214
timestamp 1644511149
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1644511149
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_244
timestamp 1644511149
transform 1 0 23552 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_253
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_260
timestamp 1644511149
transform 1 0 25024 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_400
timestamp 1644511149
transform 1 0 37904 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1644511149
transform 1 0 38456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_12
timestamp 1644511149
transform 1 0 2208 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_240
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_288
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1644511149
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 1644511149
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1644511149
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_38
timestamp 1644511149
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1644511149
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1644511149
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_228
timestamp 1644511149
transform 1 0 22080 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_250
timestamp 1644511149
transform 1 0 24104 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_262
timestamp 1644511149
transform 1 0 25208 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_354
timestamp 1644511149
transform 1 0 33672 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_379
timestamp 1644511149
transform 1 0 35972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_396
timestamp 1644511149
transform 1 0 37536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_9
timestamp 1644511149
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_173
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_212
timestamp 1644511149
transform 1 0 20608 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_216
timestamp 1644511149
transform 1 0 20976 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_222
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1644511149
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_368
timestamp 1644511149
transform 1 0 34960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_380
timestamp 1644511149
transform 1 0 36064 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_98
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1644511149
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1644511149
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1644511149
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1644511149
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_234
timestamp 1644511149
transform 1 0 22632 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_243
timestamp 1644511149
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_255
timestamp 1644511149
transform 1 0 24564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_267
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1644511149
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1644511149
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1644511149
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_88
timestamp 1644511149
transform 1 0 9200 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_115
timestamp 1644511149
transform 1 0 11684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_127
timestamp 1644511149
transform 1 0 12788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_182
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_207
timestamp 1644511149
transform 1 0 20148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_211
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_230
timestamp 1644511149
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_344
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_356
timestamp 1644511149
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_28
timestamp 1644511149
transform 1 0 3680 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_40
timestamp 1644511149
transform 1 0 4784 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1644511149
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_77
timestamp 1644511149
transform 1 0 8188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1644511149
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1644511149
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_206
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1644511149
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_240
timestamp 1644511149
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_252
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_264
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_360
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_372
timestamp 1644511149
transform 1 0 35328 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1644511149
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1644511149
transform 1 0 38456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_11
timestamp 1644511149
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1644511149
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_88
timestamp 1644511149
transform 1 0 9200 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_94
timestamp 1644511149
transform 1 0 9752 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_98
timestamp 1644511149
transform 1 0 10120 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_110
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_122
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1644511149
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1644511149
transform 1 0 21988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_342
timestamp 1644511149
transform 1 0 32568 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_354
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1644511149
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_381
timestamp 1644511149
transform 1 0 36156 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_397
timestamp 1644511149
transform 1 0 37628 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1644511149
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_37
timestamp 1644511149
transform 1 0 4508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_49
timestamp 1644511149
transform 1 0 5612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_61
timestamp 1644511149
transform 1 0 6716 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_73
timestamp 1644511149
transform 1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 1644511149
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1644511149
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_381
timestamp 1644511149
transform 1 0 36156 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_396
timestamp 1644511149
transform 1 0 37536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_36
timestamp 1644511149
transform 1 0 4416 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_48
timestamp 1644511149
transform 1 0 5520 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_60
timestamp 1644511149
transform 1 0 6624 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_72
timestamp 1644511149
transform 1 0 7728 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_371
timestamp 1644511149
transform 1 0 35236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_378
timestamp 1644511149
transform 1 0 35880 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_12
timestamp 1644511149
transform 1 0 2208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_24
timestamp 1644511149
transform 1 0 3312 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_36
timestamp 1644511149
transform 1 0 4416 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_48
timestamp 1644511149
transform 1 0 5520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1644511149
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_373
timestamp 1644511149
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_378
timestamp 1644511149
transform 1 0 35880 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1644511149
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_9
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_21
timestamp 1644511149
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_33
timestamp 1644511149
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1644511149
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1644511149
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_198
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1644511149
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_266
timestamp 1644511149
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1644511149
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_377
timestamp 1644511149
transform 1 0 35788 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_381
timestamp 1644511149
transform 1 0 36156 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1644511149
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_397
timestamp 1644511149
transform 1 0 37628 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_218
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_230
timestamp 1644511149
transform 1 0 22264 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 1644511149
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1644511149
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_259
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_271
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_283
timestamp 1644511149
transform 1 0 27140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_295
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_381
timestamp 1644511149
transform 1 0 36156 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_191
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_203
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_215
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_12
timestamp 1644511149
transform 1 0 2208 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_381
timestamp 1644511149
transform 1 0 36156 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_26
timestamp 1644511149
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_38
timestamp 1644511149
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1644511149
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_398
timestamp 1644511149
transform 1 0 37720 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1644511149
transform 1 0 38456 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_9
timestamp 1644511149
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1644511149
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_256
timestamp 1644511149
transform 1 0 24656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_268
timestamp 1644511149
transform 1 0 25760 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_280
timestamp 1644511149
transform 1 0 26864 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_292
timestamp 1644511149
transform 1 0 27968 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 1644511149
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_381
timestamp 1644511149
transform 1 0 36156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_116
timestamp 1644511149
transform 1 0 11776 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_128
timestamp 1644511149
transform 1 0 12880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_140
timestamp 1644511149
transform 1 0 13984 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_152
timestamp 1644511149
transform 1 0 15088 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_245
timestamp 1644511149
transform 1 0 23644 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_269
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1644511149
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1644511149
transform 1 0 4048 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1644511149
transform 1 0 5152 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1644511149
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1644511149
transform 1 0 7360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_120
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_127
timestamp 1644511149
transform 1 0 12788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_182
timestamp 1644511149
transform 1 0 17848 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1644511149
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_204
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_212
timestamp 1644511149
transform 1 0 20608 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_234
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_290
timestamp 1644511149
transform 1 0 27784 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_371
timestamp 1644511149
transform 1 0 35236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_378
timestamp 1644511149
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_46
timestamp 1644511149
transform 1 0 5336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_97
timestamp 1644511149
transform 1 0 10028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_101
timestamp 1644511149
transform 1 0 10396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_199
timestamp 1644511149
transform 1 0 19412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_206
timestamp 1644511149
transform 1 0 20056 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_213
timestamp 1644511149
transform 1 0 20700 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_246
timestamp 1644511149
transform 1 0 23736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_271
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1644511149
transform 1 0 30728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_356
timestamp 1644511149
transform 1 0 33856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_363
timestamp 1644511149
transform 1 0 34500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_14
timestamp 1644511149
transform 1 0 2392 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1644511149
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1644511149
transform 1 0 4048 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1644511149
transform 1 0 5152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1644511149
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1644511149
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_98
timestamp 1644511149
transform 1 0 10120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1644511149
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1644511149
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_144
timestamp 1644511149
transform 1 0 14352 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_154
timestamp 1644511149
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1644511149
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_182
timestamp 1644511149
transform 1 0 17848 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_188
timestamp 1644511149
transform 1 0 18400 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_220
timestamp 1644511149
transform 1 0 21344 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_228
timestamp 1644511149
transform 1 0 22080 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_234
timestamp 1644511149
transform 1 0 22632 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1644511149
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_256
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_268
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1644511149
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1644511149
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_397
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1644511149
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37536 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1644511149
transform 1 0 37536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1644511149
transform 1 0 37444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1644511149
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1644511149
transform -1 0 2760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1644511149
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1644511149
transform -1 0 28152 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1644511149
transform 1 0 28244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1644511149
transform -1 0 20056 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1644511149
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _293_
timestamp 1644511149
transform -1 0 20056 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1644511149
transform 1 0 33396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1644511149
transform -1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1644511149
transform -1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20608 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1644511149
transform -1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1644511149
transform -1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1644511149
transform -1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1644511149
transform -1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _305_
timestamp 1644511149
transform -1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1644511149
transform 1 0 37352 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1644511149
transform 1 0 37352 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1644511149
transform -1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _311_
timestamp 1644511149
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _312_
timestamp 1644511149
transform 1 0 18216 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1644511149
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1644511149
transform 1 0 37352 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1644511149
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1644511149
transform -1 0 4048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1644511149
transform -1 0 21344 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _318_
timestamp 1644511149
transform 1 0 19688 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1644511149
transform -1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1644511149
transform 1 0 37444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1644511149
transform -1 0 36800 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1644511149
transform -1 0 4508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _324_
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1644511149
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1644511149
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1644511149
transform 1 0 37444 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1644511149
transform -1 0 24656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1644511149
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _330_
timestamp 1644511149
transform -1 0 18768 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1644511149
transform 1 0 37444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1644511149
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1644511149
transform 1 0 37444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1644511149
transform -1 0 2208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1644511149
transform 1 0 34960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _336_
timestamp 1644511149
transform -1 0 19320 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1644511149
transform -1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform 1 0 37352 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1644511149
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _342_
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  _343_
timestamp 1644511149
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1644511149
transform -1 0 2208 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1644511149
transform 1 0 35604 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1644511149
transform -1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _349_
timestamp 1644511149
transform -1 0 19780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1644511149
transform -1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1644511149
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1644511149
transform -1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _355_
timestamp 1644511149
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1644511149
transform 1 0 37352 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1644511149
transform -1 0 19320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1644511149
transform 1 0 37444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1644511149
transform -1 0 24656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _361_
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1644511149
transform -1 0 2208 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1644511149
transform 1 0 24196 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1644511149
transform -1 0 2944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _367_
timestamp 1644511149
transform 1 0 20332 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1644511149
transform 1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _373_
timestamp 1644511149
transform -1 0 17480 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1644511149
transform -1 0 36800 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1644511149
transform -1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1644511149
transform -1 0 12788 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _379_
timestamp 1644511149
transform -1 0 18768 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1644511149
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1644511149
transform 1 0 35512 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1644511149
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1644511149
transform 1 0 34960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _385_
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1644511149
transform -1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1644511149
transform 1 0 9844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1644511149
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _391_
timestamp 1644511149
transform -1 0 18860 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1644511149
transform -1 0 17204 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1644511149
transform -1 0 32752 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1644511149
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1644511149
transform -1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1644511149
transform 1 0 20884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23276 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1644511149
transform -1 0 23184 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1644511149
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22080 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _407_
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1644511149
transform -1 0 21988 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _409_
timestamp 1644511149
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1644511149
transform -1 0 20792 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _411_
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _412_
timestamp 1644511149
transform -1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _414_
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21528 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21068 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _421_
timestamp 1644511149
transform 1 0 21528 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _423_
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _424_
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1644511149
transform -1 0 23184 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _428_
timestamp 1644511149
transform -1 0 23460 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22816 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _430_
timestamp 1644511149
transform -1 0 23552 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _431_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23460 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _433_
timestamp 1644511149
transform -1 0 25024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1644511149
transform -1 0 25300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _436_
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _437_
timestamp 1644511149
transform 1 0 23184 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_2  _439_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22816 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  _440__16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441__17
timestamp 1644511149
transform -1 0 2208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442__18
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443__19
timestamp 1644511149
transform -1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444__20
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445__21
timestamp 1644511149
transform 1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446__22
timestamp 1644511149
transform 1 0 37628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447__23
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448__24
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449__25
timestamp 1644511149
transform 1 0 35604 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450__26
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451__27
timestamp 1644511149
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _452__28
timestamp 1644511149
transform 1 0 34224 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _453__29
timestamp 1644511149
transform -1 0 4048 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _454__30
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455__31
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456__32
timestamp 1644511149
transform 1 0 37628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457__33
timestamp 1644511149
transform -1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458__34
timestamp 1644511149
transform -1 0 4416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459__35
timestamp 1644511149
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460__36
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461__37
timestamp 1644511149
transform -1 0 36800 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462__38
timestamp 1644511149
transform -1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463__39
timestamp 1644511149
transform -1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464__40
timestamp 1644511149
transform 1 0 37628 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465__41
timestamp 1644511149
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466__42
timestamp 1644511149
transform 1 0 37628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _467__43
timestamp 1644511149
transform -1 0 1932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _468__44
timestamp 1644511149
transform -1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _469__45
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470__46
timestamp 1644511149
transform -1 0 36800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471__47
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472__48
timestamp 1644511149
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473__49
timestamp 1644511149
transform -1 0 26220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474__50
timestamp 1644511149
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475__51
timestamp 1644511149
transform -1 0 1932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476__52
timestamp 1644511149
transform 1 0 37628 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477__53
timestamp 1644511149
transform -1 0 17848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478__54
timestamp 1644511149
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479__55
timestamp 1644511149
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480__56
timestamp 1644511149
transform -1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481__57
timestamp 1644511149
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482__58
timestamp 1644511149
transform -1 0 20424 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483__59
timestamp 1644511149
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484__60
timestamp 1644511149
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _485__61
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _486__62
timestamp 1644511149
transform 1 0 35880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _487__63
timestamp 1644511149
transform 1 0 18400 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _488__64
timestamp 1644511149
transform -1 0 36800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489__65
timestamp 1644511149
transform 1 0 33580 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490__66
timestamp 1644511149
transform -1 0 27876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _491__67
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492__68
timestamp 1644511149
transform -1 0 24932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _493__69
timestamp 1644511149
transform -1 0 1932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _494__70
timestamp 1644511149
transform -1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _495__71
timestamp 1644511149
transform -1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496__72
timestamp 1644511149
transform 1 0 10488 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _497__73
timestamp 1644511149
transform 1 0 37628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498__74
timestamp 1644511149
transform -1 0 36800 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _499__75
timestamp 1644511149
transform -1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500__76
timestamp 1644511149
transform -1 0 14352 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _501__77
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _502__78
timestamp 1644511149
transform -1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _503__79
timestamp 1644511149
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _504__80
timestamp 1644511149
transform -1 0 32568 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _505__81
timestamp 1644511149
transform -1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _506__82
timestamp 1644511149
transform 1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507__83
timestamp 1644511149
transform 1 0 17296 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _508__84
timestamp 1644511149
transform -1 0 20056 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509__85
timestamp 1644511149
transform -1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _510__86
timestamp 1644511149
transform -1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511__87
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512__88
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513__89
timestamp 1644511149
transform -1 0 36800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514__90
timestamp 1644511149
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515__91
timestamp 1644511149
transform 1 0 35604 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _516__92
timestamp 1644511149
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _517__93
timestamp 1644511149
transform -1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518__94
timestamp 1644511149
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _519__95
timestamp 1644511149
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520__96
timestamp 1644511149
transform -1 0 28796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _521__97
timestamp 1644511149
transform 1 0 10120 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522__98
timestamp 1644511149
transform -1 0 29808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523__99
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _524__100
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525__101
timestamp 1644511149
transform -1 0 19872 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526__102
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527__103
timestamp 1644511149
transform -1 0 36800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _528__104
timestamp 1644511149
transform 1 0 35604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529__105
timestamp 1644511149
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _530__106
timestamp 1644511149
transform -1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531__107
timestamp 1644511149
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532__108
timestamp 1644511149
transform -1 0 2116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533__109
timestamp 1644511149
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _534__110
timestamp 1644511149
transform -1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535__111
timestamp 1644511149
transform -1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _536__112
timestamp 1644511149
transform -1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _537__113
timestamp 1644511149
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538__114
timestamp 1644511149
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539__115
timestamp 1644511149
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5888 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1644511149
transform 1 0 1840 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1644511149
transform -1 0 3312 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1644511149
transform -1 0 38088 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1644511149
transform -1 0 4508 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1644511149
transform -1 0 38180 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1644511149
transform -1 0 18032 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1644511149
transform -1 0 38180 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1644511149
transform 1 0 36248 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1644511149
transform -1 0 38180 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _551_
timestamp 1644511149
transform 1 0 18952 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _552_
timestamp 1644511149
transform 1 0 36248 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _553_
timestamp 1644511149
transform 1 0 3404 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _554_
timestamp 1644511149
transform -1 0 22632 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _555_
timestamp 1644511149
transform -1 0 5244 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _556_
timestamp 1644511149
transform -1 0 38180 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _557_
timestamp 1644511149
transform 1 0 36248 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _558_
timestamp 1644511149
transform 1 0 3956 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _559_
timestamp 1644511149
transform -1 0 38180 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _560_
timestamp 1644511149
transform -1 0 9844 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _561_
timestamp 1644511149
transform 1 0 36248 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _562_
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _563_
timestamp 1644511149
transform 1 0 9200 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _564_
timestamp 1644511149
transform -1 0 38180 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _565_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _566_
timestamp 1644511149
transform -1 0 38180 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _567_
timestamp 1644511149
transform 1 0 1564 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _568_
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _569_
timestamp 1644511149
transform -1 0 6532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _570_
timestamp 1644511149
transform 1 0 36248 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _571_
timestamp 1644511149
transform 1 0 34868 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _572_
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _573_
timestamp 1644511149
transform 1 0 25852 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _574_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _575_
timestamp 1644511149
transform 1 0 1564 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _576_
timestamp 1644511149
transform -1 0 38180 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _577_
timestamp 1644511149
transform 1 0 17480 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _578_
timestamp 1644511149
transform 1 0 36248 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _579_
timestamp 1644511149
transform -1 0 3496 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _580_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _581_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _582_
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _583_
timestamp 1644511149
transform -1 0 3312 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _584_
timestamp 1644511149
transform 1 0 1564 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _585_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _586_
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _587_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _588_
timestamp 1644511149
transform 1 0 36248 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _589_
timestamp 1644511149
transform 1 0 34868 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _590_
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _591_
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _592_
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _593_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _594_
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _595_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _596_
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _597_
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _598_
timestamp 1644511149
transform 1 0 22080 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _599_
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _600_
timestamp 1644511149
transform 1 0 21344 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _601_
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _602_
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _603_
timestamp 1644511149
transform 1 0 1656 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _604_
timestamp 1644511149
transform -1 0 12144 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _605_
timestamp 1644511149
transform -1 0 38180 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _606_
timestamp 1644511149
transform 1 0 36248 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _607_
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _608_
timestamp 1644511149
transform -1 0 13708 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _609_
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _610_
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _611_
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _612_
timestamp 1644511149
transform 1 0 32292 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _613_
timestamp 1644511149
transform 1 0 19320 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _614_
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _615_
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _616_
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _617_
timestamp 1644511149
transform 1 0 9752 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _618_
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _619_
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _620_
timestamp 1644511149
transform -1 0 3772 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _621_
timestamp 1644511149
transform 1 0 36248 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _622_
timestamp 1644511149
transform 1 0 36248 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _623_
timestamp 1644511149
transform 1 0 36248 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _624_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _625_
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _626_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _627_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _628_
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _629_
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _630_
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _631_
timestamp 1644511149
transform -1 0 3312 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _632_
timestamp 1644511149
transform 1 0 3864 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _633_
timestamp 1644511149
transform 1 0 19412 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _634_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _635_
timestamp 1644511149
transform 1 0 36248 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _636_
timestamp 1644511149
transform -1 0 36800 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _637_
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _638_
timestamp 1644511149
transform 1 0 32568 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _639_
timestamp 1644511149
transform 1 0 34040 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _640_
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _641_
timestamp 1644511149
transform 1 0 32292 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _642_
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _643_
timestamp 1644511149
transform 1 0 20424 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _644_
timestamp 1644511149
transform 1 0 8464 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _645_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _646_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _647_
timestamp 1644511149
transform -1 0 3312 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform -1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform 1 0 14904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform -1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1644511149
transform -1 0 38180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1644511149
transform 1 0 35052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform -1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 6532 0 1 36992
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 36668 800 36908 6 active
port 0 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 21886 39200 21998 40000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s -10 39200 102 40000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 33268 40000 33508 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 14802 39200 14914 40000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 39200 35308 40000 35548 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 39200 3348 40000 3588 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 7718 39200 7830 40000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 9650 39200 9762 40000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 39200 12868 40000 13108 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 7074 39200 7186 40000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 5142 39200 5254 40000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 39200 8788 40000 9028 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 39274 39200 39386 40000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 39200 15588 40000 15828 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 30258 39200 30370 40000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 34766 39200 34878 40000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 39200 25108 40000 25348 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 35410 39200 35522 40000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 22530 39200 22642 40000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 39200 24428 40000 24668 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 39200 38028 40000 38268 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 39200 26468 40000 26708 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 6430 39200 6542 40000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 13548 800 13788 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 39200 22388 40000 22628 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 39200 11508 40000 11748 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 39200 10828 40000 11068 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 10938 39200 11050 40000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 39200 1988 40000 2228 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 10938 0 11050 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 28326 39200 28438 40000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 11582 39200 11694 40000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 31546 0 31658 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 39200 16948 40000 17188 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal2 s 1278 39200 1390 40000 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 19954 39200 20066 40000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 20598 39200 20710 40000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 37986 0 38098 800 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 39200 31228 40000 31468 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 23174 39200 23286 40000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 33478 0 33590 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 39200 25788 40000 26028 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 32834 39200 32946 40000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 1922 39200 2034 40000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 32834 0 32946 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 19668 800 19908 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 38630 0 38742 800 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 9006 39200 9118 40000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 17628 800 17868 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 8788 800 9028 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 19954 0 20066 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 39200 -52 40000 188 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 25788 800 26028 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 39200 14228 40000 14468 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 10294 39200 10406 40000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 8362 0 8474 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 39200 37348 40000 37588 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 39200 21708 40000 21948 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 6068 800 6308 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 32190 0 32302 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 39200 31908 40000 32148 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 33268 800 33508 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 39200 21028 40000 21268 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 36698 39200 36810 40000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 37342 0 37454 800 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 18988 800 19228 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 26394 39200 26506 40000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 32190 39200 32302 40000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 31908 800 32148 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 25106 0 25218 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 39200 18308 40000 18548 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 21886 0 21998 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 29614 39200 29726 40000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 30902 39200 31014 40000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 13514 0 13626 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 39200 628 40000 868 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 5786 0 5898 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 11508 800 11748 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 39200 5388 40000 5628 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 39200 32588 40000 32828 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 39200 30548 40000 30788 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 12226 39200 12338 40000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 39200 35988 40000 36228 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 34628 800 34868 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 39200 23748 40000 23988 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 18022 39200 18134 40000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 37986 39200 38098 40000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 14802 0 14914 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 12188 800 12428 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 39200 6068 40000 6308 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 39200 4708 40000 4948 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 12870 39200 12982 40000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 25106 39200 25218 40000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 19310 39200 19422 40000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 14158 39200 14270 40000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 38630 39200 38742 40000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 39200 7428 40000 7668 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 39200 2668 40000 2908 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 634 39200 746 40000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 33478 39200 33590 40000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 39200 19668 40000 19908 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 15446 39200 15558 40000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 16090 39200 16202 40000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 39200 9468 40000 9708 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 39200 36668 40000 36908 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal2 s 3854 39200 3966 40000 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 21242 39200 21354 40000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 39200 13548 40000 13788 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 39200 29188 40000 29428 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s 4498 39200 4610 40000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 39200 20348 40000 20588 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 35988 800 36228 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 39200 34628 40000 34868 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 24462 39200 24574 40000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 39200 14908 40000 15148 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 39200 4028 40000 4268 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 38708 800 38948 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal2 s 35410 0 35522 800 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 16734 0 16846 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 39200 10148 40000 10388 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 39200 38708 40000 38948 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal2 s 36698 0 36810 800 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 39200 16268 40000 16508 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 39200 29868 40000 30108 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 37342 39200 37454 40000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal2 s 39274 0 39386 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 36054 39200 36166 40000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 2566 39200 2678 40000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 17378 39200 17490 40000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 25750 39200 25862 40000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 16734 39200 16846 40000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 31546 39200 31658 40000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 39200 8108 40000 8348 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 39200 27828 40000 28068 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 39200 27148 40000 27388 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 27682 39200 27794 40000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 27038 39200 27150 40000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 5786 39200 5898 40000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 212 nsew ground input
rlabel metal3 s 39200 18988 40000 19228 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
